library verilog;
use verilog.vl_types.all;
entity topdct_idct is
    generic(
        BitWidth        : integer := 31
    );
end topdct_idct;
