library verilog;
use verilog.vl_types.all;
entity DLH_X2 is
    port(
        D               : in     vl_logic;
        G               : in     vl_logic;
        Q               : out    vl_logic
    );
end DLH_X2;
