module conf_int_mul__noFF__arch_agnos_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 ( clk, 
        rst, a, b, \d[47] , \d[44] , \d[43] , \d[40] , \d[37]_BAR , \d[34] , 
        \d[31] , \d[28] , \d[16] , \d[1] , \d[0] , \d[33]_BAR , \d[27]_BAR , 
        \d[26]_BAR , \d[24]_BAR , \d[23]_BAR , \d[15]_BAR , \d[14]_BAR , 
        \d[11]_BAR , \d[9]_BAR , \d[6]_BAR , \d[4]_BAR , \d[42]_BAR , 
        \d[41]_BAR , \d[30] , \d[22]_BAR , \d[46]_BAR , \d[35] , \d[19] , 
        \d[8]_BAR , \d[5]_BAR , \d[3] , \d[29] , \d[32] , \d[39]_BAR , \d[2] , 
        \d[36]_BAR , \d[25] , \d[13]_BAR , \d[38]_BAR , \d[20] , \d[18] , 
        \d[17]_BAR , \d[45]_BAR , \d[21] , \d[12] , \d[10] , \d[7]  );
  input [23:0] a;
  input [23:0] b;
  input clk, rst;
  output \d[47] , \d[44] , \d[43] , \d[40] , \d[37]_BAR , \d[34] , \d[31] ,
         \d[28] , \d[16] , \d[1] , \d[0] , \d[33]_BAR , \d[27]_BAR ,
         \d[26]_BAR , \d[24]_BAR , \d[23]_BAR , \d[15]_BAR , \d[14]_BAR ,
         \d[11]_BAR , \d[9]_BAR , \d[6]_BAR , \d[4]_BAR , \d[42]_BAR ,
         \d[41]_BAR , \d[30] , \d[22]_BAR , \d[46]_BAR , \d[35] , \d[19] ,
         \d[8]_BAR , \d[5]_BAR , \d[3] , \d[29] , \d[32] , \d[39]_BAR , \d[2] ,
         \d[36]_BAR , \d[25] , \d[13]_BAR , \d[38]_BAR , \d[20] , \d[18] ,
         \d[17]_BAR , \d[45]_BAR , \d[21] , \d[12] , \d[10] , \d[7] ;
  wire   \intadd_46/A[4] , \intadd_46/A[3] , \intadd_46/A[2] ,
         \intadd_46/A[1] , \intadd_46/A[0] , \intadd_46/B[3] ,
         \intadd_46/B[2] , \intadd_46/B[1] , \intadd_46/B[0] , \intadd_46/CI ,
         \intadd_46/SUM[2] , \intadd_46/SUM[1] , \intadd_46/SUM[0] ,
         \intadd_46/n5 , \intadd_46/n4 , \intadd_46/n3 , \intadd_46/n2 ,
         \intadd_47/A[4] , \intadd_47/A[3] , \intadd_47/A[2] ,
         \intadd_47/A[1] , \intadd_47/B[4] , \intadd_47/B[3] ,
         \intadd_47/B[2] , \intadd_47/B[1] , \intadd_47/B[0] , \intadd_47/CI ,
         \intadd_47/SUM[4] , \intadd_47/SUM[3] , \intadd_47/SUM[2] ,
         \intadd_47/SUM[1] , \intadd_47/SUM[0] , \intadd_47/n5 ,
         \intadd_47/n4 , \intadd_47/n3 , \intadd_47/n2 , \intadd_47/n1 ,
         \intadd_48/A[4] , \intadd_48/A[3] , \intadd_48/A[2] ,
         \intadd_48/A[1] , \intadd_48/A[0] , \intadd_48/B[4] ,
         \intadd_48/B[3] , \intadd_48/B[2] , \intadd_48/B[1] ,
         \intadd_48/B[0] , \intadd_48/SUM[4] , \intadd_48/SUM[2] ,
         \intadd_48/SUM[0] , \intadd_48/n5 , \intadd_48/n4 , \intadd_48/n3 ,
         \intadd_48/n2 , \intadd_48/n1 , \intadd_49/A[3] , \intadd_49/A[2] ,
         \intadd_49/A[1] , \intadd_49/B[0] , \intadd_49/CI ,
         \intadd_49/SUM[4] , \intadd_49/SUM[3] , \intadd_49/SUM[2] ,
         \intadd_49/SUM[1] , \intadd_49/SUM[0] , \intadd_49/n5 ,
         \intadd_49/n4 , \intadd_49/n3 , \intadd_49/n2 , \intadd_49/n1 ,
         \intadd_50/A[1] , \intadd_50/A[0] , \intadd_50/B[3] ,
         \intadd_50/B[2] , \intadd_50/B[1] , \intadd_50/CI ,
         \intadd_50/SUM[4] , \intadd_50/SUM[3] , \intadd_50/SUM[2] ,
         \intadd_50/SUM[1] , \intadd_50/SUM[0] , \intadd_50/n5 ,
         \intadd_50/n4 , \intadd_50/n3 , \intadd_50/n2 , \intadd_50/n1 ,
         \intadd_51/A[4] , \intadd_51/A[3] , \intadd_51/A[2] ,
         \intadd_51/A[1] , \intadd_51/A[0] , \intadd_51/B[4] ,
         \intadd_51/B[3] , \intadd_51/B[2] , \intadd_51/B[1] , \intadd_51/CI ,
         \intadd_51/SUM[4] , \intadd_51/SUM[3] , \intadd_51/SUM[2] ,
         \intadd_51/SUM[1] , \intadd_51/SUM[0] , \intadd_51/n5 ,
         \intadd_51/n4 , \intadd_51/n3 , \intadd_51/n2 , \intadd_51/n1 ,
         \intadd_52/A[4] , \intadd_52/A[2] , \intadd_52/A[1] ,
         \intadd_52/A[0] , \intadd_52/B[4] , \intadd_52/B[3] ,
         \intadd_52/B[2] , \intadd_52/B[1] , \intadd_52/B[0] ,
         \intadd_52/SUM[4] , \intadd_52/SUM[3] , \intadd_52/SUM[2] ,
         \intadd_52/SUM[1] , \intadd_52/SUM[0] , \intadd_52/n5 ,
         \intadd_52/n4 , \intadd_52/n3 , \intadd_52/n2 , \intadd_52/n1 ,
         \intadd_53/A[4] , \intadd_53/A[3] , \intadd_53/A[2] ,
         \intadd_53/A[1] , \intadd_53/A[0] , \intadd_53/B[3] ,
         \intadd_53/B[2] , \intadd_53/B[1] , \intadd_53/B[0] , \intadd_53/CI ,
         \intadd_53/SUM[4] , \intadd_53/SUM[3] , \intadd_53/SUM[2] ,
         \intadd_53/SUM[1] , \intadd_53/SUM[0] , \intadd_53/n5 ,
         \intadd_53/n4 , \intadd_53/n3 , \intadd_53/n2 , \intadd_53/n1 ,
         \intadd_54/A[4] , \intadd_54/A[2] , \intadd_54/A[1] ,
         \intadd_54/A[0] , \intadd_54/B[4] , \intadd_54/B[2] ,
         \intadd_54/B[1] , \intadd_54/B[0] , \intadd_54/CI ,
         \intadd_54/SUM[4] , \intadd_54/SUM[2] , \intadd_54/SUM[1] ,
         \intadd_54/SUM[0] , \intadd_54/n5 , \intadd_54/n4 , \intadd_54/n3 ,
         \intadd_54/n2 , \intadd_54/n1 , \intadd_55/A[4] , \intadd_55/A[3] ,
         \intadd_55/A[2] , \intadd_55/A[1] , \intadd_55/A[0] ,
         \intadd_55/B[4] , \intadd_55/B[3] , \intadd_55/B[2] ,
         \intadd_55/B[1] , \intadd_55/B[0] , \intadd_55/CI ,
         \intadd_55/SUM[4] , \intadd_55/SUM[3] , \intadd_55/SUM[2] ,
         \intadd_55/SUM[1] , \intadd_55/SUM[0] , \intadd_55/n5 ,
         \intadd_55/n4 , \intadd_55/n3 , \intadd_55/n2 , \intadd_55/n1 ,
         \intadd_56/A[4] , \intadd_56/A[3] , \intadd_56/A[2] ,
         \intadd_56/A[1] , \intadd_56/A[0] , \intadd_56/B[4] ,
         \intadd_56/B[3] , \intadd_56/B[2] , \intadd_56/B[1] , \intadd_56/CI ,
         \intadd_56/SUM[4] , \intadd_56/SUM[2] , \intadd_56/SUM[1] ,
         \intadd_56/n5 , \intadd_56/n4 , \intadd_56/n3 , \intadd_56/n2 ,
         \intadd_56/n1 , \intadd_57/A[1] , \intadd_57/B[3] , \intadd_57/B[0] ,
         \intadd_57/CI , \intadd_57/SUM[1] , \intadd_57/SUM[0] ,
         \intadd_57/n4 , \intadd_57/n3 , \intadd_57/n2 , \intadd_57/n1 ,
         \intadd_58/A[3] , \intadd_58/A[2] , \intadd_58/A[1] ,
         \intadd_58/B[3] , \intadd_58/B[2] , \intadd_58/B[1] ,
         \intadd_58/B[0] , \intadd_58/CI , \intadd_58/SUM[3] ,
         \intadd_58/SUM[2] , \intadd_58/SUM[1] , \intadd_58/SUM[0] ,
         \intadd_58/n4 , \intadd_58/n3 , \intadd_58/n2 , \intadd_58/n1 ,
         \intadd_59/A[3] , \intadd_59/A[2] , \intadd_59/A[1] ,
         \intadd_59/A[0] , \intadd_59/B[3] , \intadd_59/B[2] ,
         \intadd_59/B[1] , \intadd_59/B[0] , \intadd_59/SUM[3] ,
         \intadd_59/SUM[0] , \intadd_59/n4 , \intadd_59/n3 , \intadd_59/n2 ,
         \intadd_59/n1 , \intadd_60/A[3] , \intadd_60/A[2] , \intadd_60/A[1] ,
         \intadd_60/B[3] , \intadd_60/B[2] , \intadd_60/B[1] ,
         \intadd_60/B[0] , \intadd_60/SUM[3] , \intadd_60/SUM[0] ,
         \intadd_60/n4 , \intadd_60/n3 , \intadd_60/n2 , \intadd_60/n1 ,
         \intadd_61/A[3] , \intadd_61/A[2] , \intadd_61/A[1] ,
         \intadd_61/A[0] , \intadd_61/B[3] , \intadd_61/B[2] ,
         \intadd_61/B[1] , \intadd_61/CI , \intadd_61/SUM[0] , \intadd_61/n4 ,
         \intadd_61/n3 , \intadd_61/n2 , \intadd_61/n1 , \intadd_62/A[3] ,
         \intadd_62/A[2] , \intadd_62/A[1] , \intadd_62/A[0] ,
         \intadd_62/B[3] , \intadd_62/B[2] , \intadd_62/B[1] ,
         \intadd_62/B[0] , \intadd_62/n4 , \intadd_62/n3 , \intadd_62/n2 ,
         \intadd_62/n1 , \intadd_63/A[1] , \intadd_63/A[0] , \intadd_63/B[3] ,
         \intadd_63/B[2] , \intadd_63/B[1] , \intadd_63/B[0] , \intadd_63/CI ,
         \intadd_63/SUM[3] , \intadd_63/SUM[1] , \intadd_63/SUM[0] ,
         \intadd_63/n4 , \intadd_63/n3 , \intadd_63/n2 , \intadd_63/n1 ,
         \intadd_64/A[3] , \intadd_64/A[2] , \intadd_64/A[1] ,
         \intadd_64/A[0] , \intadd_64/B[3] , \intadd_64/B[2] ,
         \intadd_64/B[1] , \intadd_64/B[0] , \intadd_64/CI ,
         \intadd_64/SUM[2] , \intadd_64/n4 , \intadd_64/n3 , \intadd_64/n2 ,
         \intadd_64/n1 , \intadd_65/A[3] , \intadd_65/A[2] , \intadd_65/A[1] ,
         \intadd_65/A[0] , \intadd_65/B[3] , \intadd_65/B[2] ,
         \intadd_65/B[1] , \intadd_65/B[0] , \intadd_65/CI ,
         \intadd_65/SUM[3] , \intadd_65/SUM[2] , \intadd_65/SUM[1] ,
         \intadd_65/SUM[0] , \intadd_65/n4 , \intadd_65/n3 , \intadd_65/n2 ,
         \intadd_65/n1 , \intadd_66/A[3] , \intadd_66/A[2] , \intadd_66/A[1] ,
         \intadd_66/A[0] , \intadd_66/B[2] , \intadd_66/B[1] ,
         \intadd_66/B[0] , \intadd_66/CI , \intadd_66/SUM[3] ,
         \intadd_66/SUM[2] , \intadd_66/n4 , \intadd_66/n3 , \intadd_66/n2 ,
         \intadd_66/n1 , \intadd_67/A[3] , \intadd_67/A[2] , \intadd_67/A[1] ,
         \intadd_67/A[0] , \intadd_67/B[2] , \intadd_67/B[1] ,
         \intadd_67/B[0] , \intadd_67/CI , \intadd_67/SUM[3] ,
         \intadd_67/SUM[2] , \intadd_67/SUM[1] , \intadd_67/SUM[0] ,
         \intadd_67/n4 , \intadd_67/n3 , \intadd_67/n2 , \intadd_67/n1 ,
         \intadd_68/A[3] , \intadd_68/A[2] , \intadd_68/A[1] ,
         \intadd_68/A[0] , \intadd_68/B[3] , \intadd_68/B[2] ,
         \intadd_68/B[1] , \intadd_68/CI , \intadd_68/SUM[3] ,
         \intadd_68/SUM[2] , \intadd_68/SUM[1] , \intadd_68/SUM[0] ,
         \intadd_68/n4 , \intadd_68/n3 , \intadd_68/n2 , \intadd_68/n1 ,
         \intadd_69/A[3] , \intadd_69/A[2] , \intadd_69/A[1] ,
         \intadd_69/A[0] , \intadd_69/B[2] , \intadd_69/B[1] , \intadd_69/CI ,
         \intadd_69/SUM[3] , \intadd_69/SUM[2] , \intadd_69/SUM[1] ,
         \intadd_69/SUM[0] , \intadd_69/n4 , \intadd_69/n3 , \intadd_69/n2 ,
         \intadd_69/n1 , \intadd_70/A[2] , \intadd_70/A[1] , \intadd_70/A[0] ,
         \intadd_70/B[2] , \intadd_70/B[1] , \intadd_70/B[0] , \intadd_70/CI ,
         \intadd_70/n3 , \intadd_70/n2 , \intadd_70/n1 , \intadd_71/A[1] ,
         \intadd_71/A[0] , \intadd_71/B[2] , \intadd_71/B[1] , \intadd_71/CI ,
         \intadd_71/SUM[2] , \intadd_71/SUM[1] , \intadd_71/SUM[0] ,
         \intadd_71/n3 , \intadd_71/n2 , \intadd_71/n1 , \intadd_72/A[2] ,
         \intadd_72/A[0] , \intadd_72/B[2] , \intadd_72/B[0] , \intadd_72/CI ,
         \intadd_72/SUM[2] , \intadd_72/SUM[0] , \intadd_72/n3 ,
         \intadd_72/n2 , \intadd_72/n1 , \intadd_73/A[1] , \intadd_73/A[0] ,
         \intadd_73/B[2] , \intadd_73/B[1] , \intadd_73/B[0] , \intadd_73/CI ,
         \intadd_73/SUM[1] , \intadd_73/SUM[0] , \intadd_73/n3 ,
         \intadd_73/n2 , \intadd_73/n1 , \intadd_74/A[2] , \intadd_74/A[1] ,
         \intadd_74/A[0] , \intadd_74/B[2] , \intadd_74/B[1] ,
         \intadd_74/B[0] , \intadd_74/CI , \intadd_74/SUM[2] ,
         \intadd_74/SUM[1] , \intadd_74/SUM[0] , \intadd_74/n3 ,
         \intadd_74/n2 , \intadd_74/n1 , \intadd_75/A[2] , \intadd_75/A[1] ,
         \intadd_75/A[0] , \intadd_75/B[1] , \intadd_75/B[0] , \intadd_75/CI ,
         \intadd_75/SUM[1] , \intadd_75/SUM[0] , \intadd_75/n3 ,
         \intadd_75/n2 , \intadd_75/n1 , \intadd_76/A[2] , \intadd_76/A[1] ,
         \intadd_76/A[0] , \intadd_76/B[2] , \intadd_76/B[1] ,
         \intadd_76/B[0] , \intadd_76/CI , \intadd_76/SUM[2] ,
         \intadd_76/SUM[1] , \intadd_76/SUM[0] , \intadd_76/n3 ,
         \intadd_76/n2 , \intadd_76/n1 , \intadd_77/A[1] , \intadd_77/A[0] ,
         \intadd_77/B[0] , \intadd_77/SUM[2] , \intadd_77/SUM[1] ,
         \intadd_77/n3 , \intadd_77/n2 , \intadd_77/n1 , \intadd_78/A[2] ,
         \intadd_78/A[1] , \intadd_78/A[0] , \intadd_78/B[2] ,
         \intadd_78/B[1] , \intadd_78/B[0] , \intadd_78/CI ,
         \intadd_78/SUM[2] , \intadd_78/SUM[1] , \intadd_78/SUM[0] ,
         \intadd_78/n3 , \intadd_78/n2 , \intadd_78/n1 , \intadd_79/A[2] ,
         \intadd_79/A[0] , \intadd_79/B[2] , \intadd_79/B[1] ,
         \intadd_79/B[0] , \intadd_79/CI , \intadd_79/SUM[0] , \intadd_79/n3 ,
         \intadd_79/n2 , \intadd_79/n1 , \intadd_80/A[2] , \intadd_80/A[1] ,
         \intadd_80/A[0] , \intadd_80/B[2] , \intadd_80/B[1] ,
         \intadd_80/B[0] , \intadd_80/CI , \intadd_80/n3 , \intadd_80/n2 ,
         \intadd_80/n1 , \intadd_81/A[0] , \intadd_81/B[2] , \intadd_81/B[1] ,
         \intadd_81/B[0] , \intadd_81/CI , \intadd_81/SUM[2] ,
         \intadd_81/SUM[0] , \intadd_81/n3 , \intadd_81/n2 , \intadd_81/n1 ,
         n2, n4, n5, n8, n9, n10, n11, n12, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n31, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n90, n91, n92, n93, n96, n97, n98, n101, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n162, n163, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n177, n178, n179, n180, n181,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n215, n216,
         n217, n218, n219, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n312, n314, n315, n316, n317, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n338, n339, n340, n341, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n518,
         n519, n520, n521, n522, n523, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n569, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n735, n736, n737, n738, n739, n740, n741,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1627, n1628, n1629, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2083, n2084, n2085, n2086, n2087, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255;
  assign \d[12]  = \intadd_54/SUM[4] ;
  assign \d[10]  = \intadd_54/SUM[2] ;
  assign \d[45]_BAR  = \intadd_58/SUM[3] ;
  assign \d[7]  = \intadd_72/SUM[2] ;

  FA_X1 \intadd_46/U6  ( .A(\intadd_46/A[0] ), .B(\intadd_46/B[0] ), .CI(
        \intadd_46/CI ), .CO(\intadd_46/n5 ), .S(\intadd_46/SUM[0] ) );
  FA_X1 \intadd_46/U5  ( .A(\intadd_46/A[1] ), .B(\intadd_46/B[1] ), .CI(
        \intadd_46/n5 ), .CO(\intadd_46/n4 ), .S(\intadd_46/SUM[1] ) );
  FA_X1 \intadd_46/U4  ( .A(\intadd_46/A[2] ), .B(\intadd_46/B[2] ), .CI(
        \intadd_46/n4 ), .CO(\intadd_46/n3 ), .S(\intadd_46/SUM[2] ) );
  FA_X1 \intadd_46/U3  ( .A(\intadd_46/A[3] ), .B(\intadd_46/B[3] ), .CI(
        \intadd_46/n3 ), .CO(\intadd_46/n2 ), .S(\d[13]_BAR ) );
  FA_X1 \intadd_47/U6  ( .A(n2192), .B(\intadd_47/B[0] ), .CI(\intadd_47/CI ), 
        .CO(\intadd_47/n5 ), .S(\intadd_47/SUM[0] ) );
  FA_X1 \intadd_47/U5  ( .A(\intadd_47/A[1] ), .B(\intadd_47/B[1] ), .CI(
        \intadd_47/n5 ), .CO(\intadd_47/n4 ), .S(\intadd_47/SUM[1] ) );
  FA_X1 \intadd_47/U4  ( .A(\intadd_47/A[2] ), .B(\intadd_47/B[2] ), .CI(
        \intadd_47/n4 ), .CO(\intadd_47/n3 ), .S(\intadd_47/SUM[2] ) );
  FA_X1 \intadd_47/U3  ( .A(\intadd_47/A[3] ), .B(\intadd_47/B[3] ), .CI(
        \intadd_47/n3 ), .CO(\intadd_47/n2 ), .S(\intadd_47/SUM[3] ) );
  FA_X1 \intadd_47/U2  ( .A(\intadd_47/A[4] ), .B(\intadd_47/B[4] ), .CI(
        \intadd_47/n2 ), .CO(\intadd_47/n1 ), .S(\intadd_47/SUM[4] ) );
  FA_X1 \intadd_48/U6  ( .A(\intadd_48/A[0] ), .B(\intadd_48/B[0] ), .CI(n2194), .CO(\intadd_48/n5 ), .S(\intadd_48/SUM[0] ) );
  FA_X1 \intadd_48/U5  ( .A(\intadd_48/A[1] ), .B(\intadd_48/B[1] ), .CI(
        \intadd_48/n5 ), .CO(\intadd_48/n4 ), .S(\intadd_47/A[2] ) );
  FA_X1 \intadd_48/U4  ( .A(\intadd_48/A[2] ), .B(\intadd_48/B[2] ), .CI(
        \intadd_48/n4 ), .CO(\intadd_48/n3 ), .S(\intadd_48/SUM[2] ) );
  FA_X1 \intadd_48/U3  ( .A(\intadd_48/A[3] ), .B(\intadd_48/B[3] ), .CI(
        \intadd_48/n3 ), .CO(\intadd_48/n2 ), .S(\intadd_47/A[4] ) );
  FA_X1 \intadd_48/U2  ( .A(\intadd_48/A[4] ), .B(\intadd_48/B[4] ), .CI(
        \intadd_48/n2 ), .CO(\intadd_48/n1 ), .S(\intadd_48/SUM[4] ) );
  FA_X1 \intadd_49/U6  ( .A(n2193), .B(\intadd_49/B[0] ), .CI(\intadd_49/CI ), 
        .CO(\intadd_49/n5 ), .S(\intadd_49/SUM[0] ) );
  FA_X1 \intadd_49/U5  ( .A(\intadd_49/A[1] ), .B(n2190), .CI(\intadd_49/n5 ), 
        .CO(\intadd_49/n4 ), .S(\intadd_49/SUM[1] ) );
  FA_X1 \intadd_49/U4  ( .A(\intadd_49/A[2] ), .B(\intadd_48/SUM[0] ), .CI(
        \intadd_49/n4 ), .CO(\intadd_49/n3 ), .S(\intadd_49/SUM[2] ) );
  FA_X1 \intadd_49/U3  ( .A(\intadd_49/A[3] ), .B(\intadd_71/n1 ), .CI(
        \intadd_49/n3 ), .CO(\intadd_49/n2 ), .S(\intadd_49/SUM[3] ) );
  FA_X1 \intadd_49/U2  ( .A(\intadd_47/SUM[3] ), .B(\intadd_48/SUM[2] ), .CI(
        \intadd_49/n2 ), .CO(\intadd_49/n1 ), .S(\intadd_49/SUM[4] ) );
  FA_X1 \intadd_50/U6  ( .A(\intadd_50/A[0] ), .B(n2185), .CI(\intadd_50/CI ), 
        .CO(\intadd_50/n5 ), .S(\intadd_50/SUM[0] ) );
  FA_X1 \intadd_50/U5  ( .A(\intadd_50/A[1] ), .B(\intadd_50/B[1] ), .CI(
        \intadd_50/n5 ), .CO(\intadd_50/n4 ), .S(\intadd_50/SUM[1] ) );
  FA_X1 \intadd_50/U4  ( .A(\intadd_47/SUM[0] ), .B(\intadd_50/B[2] ), .CI(
        \intadd_50/n4 ), .CO(\intadd_50/n3 ), .S(\intadd_50/SUM[2] ) );
  FA_X1 \intadd_50/U3  ( .A(\intadd_49/SUM[2] ), .B(\intadd_50/B[3] ), .CI(
        \intadd_50/n3 ), .CO(\intadd_50/n2 ), .S(\intadd_50/SUM[3] ) );
  FA_X1 \intadd_50/U2  ( .A(\intadd_47/SUM[2] ), .B(\intadd_49/SUM[3] ), .CI(
        \intadd_50/n2 ), .CO(\intadd_50/n1 ), .S(\intadd_50/SUM[4] ) );
  FA_X1 \intadd_51/U6  ( .A(\intadd_51/A[0] ), .B(n2184), .CI(\intadd_51/CI ), 
        .CO(\intadd_51/n5 ), .S(\intadd_51/SUM[0] ) );
  FA_X1 \intadd_51/U5  ( .A(\intadd_51/A[1] ), .B(\intadd_51/B[1] ), .CI(
        \intadd_51/n5 ), .CO(\intadd_51/n4 ), .S(\intadd_51/SUM[1] ) );
  FA_X1 \intadd_51/U4  ( .A(\intadd_51/A[2] ), .B(\intadd_51/B[2] ), .CI(
        \intadd_51/n4 ), .CO(\intadd_51/n3 ), .S(\intadd_51/SUM[2] ) );
  FA_X1 \intadd_51/U3  ( .A(\intadd_51/A[3] ), .B(\intadd_51/B[3] ), .CI(
        \intadd_51/n3 ), .CO(\intadd_51/n2 ), .S(\intadd_51/SUM[3] ) );
  FA_X1 \intadd_51/U2  ( .A(\intadd_51/A[4] ), .B(\intadd_51/B[4] ), .CI(
        \intadd_51/n2 ), .CO(\intadd_51/n1 ), .S(\intadd_51/SUM[4] ) );
  FA_X1 \intadd_52/U6  ( .A(\intadd_52/A[0] ), .B(\intadd_52/B[0] ), .CI(n2198), .CO(\intadd_52/n5 ), .S(\intadd_52/SUM[0] ) );
  FA_X1 \intadd_52/U5  ( .A(\intadd_52/A[1] ), .B(\intadd_52/B[1] ), .CI(
        \intadd_52/n5 ), .CO(\intadd_52/n4 ), .S(\intadd_52/SUM[1] ) );
  FA_X1 \intadd_52/U4  ( .A(\intadd_52/A[2] ), .B(\intadd_52/B[2] ), .CI(
        \intadd_52/n4 ), .CO(\intadd_52/n3 ), .S(\intadd_52/SUM[2] ) );
  FA_X1 \intadd_52/U3  ( .A(\intadd_70/n1 ), .B(\intadd_52/B[3] ), .CI(
        \intadd_52/n3 ), .CO(\intadd_52/n2 ), .S(\intadd_52/SUM[3] ) );
  FA_X1 \intadd_52/U2  ( .A(\intadd_52/A[4] ), .B(\intadd_52/B[4] ), .CI(
        \intadd_52/n2 ), .CO(\intadd_52/n1 ), .S(\intadd_52/SUM[4] ) );
  FA_X1 \intadd_53/U6  ( .A(\intadd_53/A[0] ), .B(\intadd_53/B[0] ), .CI(
        \intadd_53/CI ), .CO(\intadd_53/n5 ), .S(\intadd_53/SUM[0] ) );
  FA_X1 \intadd_53/U5  ( .A(\intadd_53/A[1] ), .B(\intadd_53/B[1] ), .CI(
        \intadd_53/n5 ), .CO(\intadd_53/n4 ), .S(\intadd_53/SUM[1] ) );
  FA_X1 \intadd_53/U4  ( .A(\intadd_53/A[2] ), .B(\intadd_53/B[2] ), .CI(
        \intadd_53/n4 ), .CO(\intadd_53/n3 ), .S(\intadd_53/SUM[2] ) );
  FA_X1 \intadd_53/U3  ( .A(\intadd_53/A[3] ), .B(\intadd_53/B[3] ), .CI(
        \intadd_53/n3 ), .CO(\intadd_53/n2 ), .S(\intadd_53/SUM[3] ) );
  FA_X1 \intadd_53/U2  ( .A(\intadd_53/A[4] ), .B(\intadd_52/SUM[3] ), .CI(
        \intadd_53/n2 ), .CO(\intadd_53/n1 ), .S(\intadd_53/SUM[4] ) );
  FA_X1 \intadd_54/U6  ( .A(\intadd_54/A[0] ), .B(\intadd_54/B[0] ), .CI(
        \intadd_54/CI ), .CO(\intadd_54/n5 ), .S(\intadd_54/SUM[0] ) );
  FA_X1 \intadd_54/U5  ( .A(\intadd_54/A[1] ), .B(\intadd_54/B[1] ), .CI(
        \intadd_54/n5 ), .CO(\intadd_54/n4 ), .S(\intadd_54/SUM[1] ) );
  FA_X1 \intadd_54/U4  ( .A(\intadd_54/A[2] ), .B(\intadd_54/B[2] ), .CI(
        \intadd_54/n4 ), .CO(\intadd_54/n3 ), .S(\intadd_54/SUM[2] ) );
  FA_X1 \intadd_54/U2  ( .A(\intadd_54/A[4] ), .B(\intadd_54/B[4] ), .CI(
        \intadd_54/n2 ), .CO(\intadd_54/n1 ), .S(\intadd_54/SUM[4] ) );
  FA_X1 \intadd_55/U6  ( .A(\intadd_55/A[0] ), .B(\intadd_55/B[0] ), .CI(
        \intadd_55/CI ), .CO(\intadd_55/n5 ), .S(\intadd_55/SUM[0] ) );
  FA_X1 \intadd_55/U5  ( .A(\intadd_55/A[1] ), .B(\intadd_55/B[1] ), .CI(
        \intadd_55/n5 ), .CO(\intadd_55/n4 ), .S(\intadd_55/SUM[1] ) );
  FA_X1 \intadd_55/U4  ( .A(\intadd_55/A[2] ), .B(\intadd_55/B[2] ), .CI(
        \intadd_55/n4 ), .CO(\intadd_55/n3 ), .S(\intadd_55/SUM[2] ) );
  FA_X1 \intadd_55/U3  ( .A(\intadd_55/A[3] ), .B(\intadd_55/B[3] ), .CI(
        \intadd_55/n3 ), .CO(\intadd_55/n2 ), .S(\intadd_55/SUM[3] ) );
  FA_X1 \intadd_55/U2  ( .A(\intadd_55/A[4] ), .B(\intadd_55/B[4] ), .CI(
        \intadd_55/n2 ), .CO(\intadd_55/n1 ), .S(\intadd_55/SUM[4] ) );
  FA_X1 \intadd_56/U6  ( .A(\intadd_56/A[0] ), .B(n2189), .CI(\intadd_56/CI ), 
        .CO(\intadd_56/n5 ), .S(\intadd_55/A[1] ) );
  FA_X1 \intadd_56/U5  ( .A(\intadd_56/A[1] ), .B(\intadd_56/B[1] ), .CI(
        \intadd_56/n5 ), .CO(\intadd_56/n4 ), .S(\intadd_56/SUM[1] ) );
  FA_X1 \intadd_56/U4  ( .A(\intadd_56/A[2] ), .B(\intadd_56/B[2] ), .CI(
        \intadd_56/n4 ), .CO(\intadd_56/n3 ), .S(\intadd_56/SUM[2] ) );
  FA_X1 \intadd_56/U3  ( .A(\intadd_56/A[3] ), .B(\intadd_56/B[3] ), .CI(
        \intadd_56/n3 ), .CO(\intadd_56/n2 ), .S(\intadd_55/A[4] ) );
  FA_X1 \intadd_56/U2  ( .A(\intadd_56/A[4] ), .B(\intadd_56/B[4] ), .CI(
        \intadd_56/n2 ), .CO(\intadd_56/n1 ), .S(\intadd_56/SUM[4] ) );
  FA_X1 \intadd_57/U5  ( .A(\intadd_77/n1 ), .B(\intadd_57/B[0] ), .CI(
        \intadd_57/CI ), .CO(\intadd_57/n4 ), .S(\intadd_57/SUM[0] ) );
  FA_X1 \intadd_57/U4  ( .A(\intadd_57/A[1] ), .B(\intadd_55/SUM[4] ), .CI(
        \intadd_57/n4 ), .CO(\intadd_57/n3 ), .S(\intadd_57/SUM[1] ) );
  FA_X1 \intadd_57/U3  ( .A(\intadd_55/n1 ), .B(\intadd_56/SUM[4] ), .CI(
        \intadd_57/n3 ), .CO(\intadd_57/n2 ), .S(\d[22]_BAR ) );
  FA_X1 \intadd_57/U2  ( .A(\intadd_56/n1 ), .B(\intadd_57/B[3] ), .CI(
        \intadd_57/n2 ), .CO(\intadd_57/n1 ), .S(\d[23]_BAR ) );
  FA_X1 \intadd_58/U5  ( .A(n2191), .B(\intadd_58/B[0] ), .CI(\intadd_58/CI ), 
        .CO(\intadd_58/n4 ), .S(\intadd_58/SUM[0] ) );
  FA_X1 \intadd_58/U4  ( .A(\intadd_58/A[1] ), .B(\intadd_58/B[1] ), .CI(
        \intadd_58/n4 ), .CO(\intadd_58/n3 ), .S(\intadd_58/SUM[1] ) );
  FA_X1 \intadd_58/U3  ( .A(\intadd_58/A[2] ), .B(\intadd_58/B[2] ), .CI(
        \intadd_58/n3 ), .CO(\intadd_58/n2 ), .S(\intadd_58/SUM[2] ) );
  FA_X1 \intadd_58/U2  ( .A(\intadd_58/A[3] ), .B(\intadd_58/B[3] ), .CI(
        \intadd_58/n2 ), .CO(\intadd_58/n1 ), .S(\intadd_58/SUM[3] ) );
  FA_X1 \intadd_59/U5  ( .A(\intadd_59/A[0] ), .B(\intadd_59/B[0] ), .CI(n2195), .CO(\intadd_59/n4 ), .S(\intadd_59/SUM[0] ) );
  FA_X1 \intadd_59/U4  ( .A(\intadd_59/A[1] ), .B(\intadd_59/B[1] ), .CI(
        \intadd_59/n4 ), .CO(\intadd_59/n3 ), .S(\intadd_48/A[3] ) );
  FA_X1 \intadd_59/U3  ( .A(\intadd_59/A[2] ), .B(\intadd_59/B[2] ), .CI(
        \intadd_59/n3 ), .CO(\intadd_59/n2 ), .S(\intadd_48/A[4] ) );
  FA_X1 \intadd_59/U2  ( .A(\intadd_59/A[3] ), .B(\intadd_59/B[3] ), .CI(
        \intadd_59/n2 ), .CO(\intadd_59/n1 ), .S(\intadd_59/SUM[3] ) );
  FA_X1 \intadd_60/U5  ( .A(n2182), .B(\intadd_60/B[0] ), .CI(n2197), .CO(
        \intadd_60/n4 ), .S(\intadd_60/SUM[0] ) );
  FA_X1 \intadd_60/U4  ( .A(\intadd_60/A[1] ), .B(\intadd_60/B[1] ), .CI(
        \intadd_60/n4 ), .CO(\intadd_60/n3 ), .S(\intadd_59/B[2] ) );
  FA_X1 \intadd_60/U3  ( .A(\intadd_60/A[2] ), .B(\intadd_60/B[2] ), .CI(
        \intadd_60/n3 ), .CO(\intadd_60/n2 ), .S(\intadd_59/A[3] ) );
  FA_X1 \intadd_60/U2  ( .A(\intadd_60/A[3] ), .B(\intadd_60/B[3] ), .CI(
        \intadd_60/n2 ), .CO(\intadd_60/n1 ), .S(\intadd_60/SUM[3] ) );
  FA_X1 \intadd_61/U5  ( .A(\intadd_61/A[0] ), .B(n2186), .CI(\intadd_61/CI ), 
        .CO(\intadd_61/n4 ), .S(\intadd_61/SUM[0] ) );
  FA_X1 \intadd_61/U4  ( .A(\intadd_61/A[1] ), .B(\intadd_61/B[1] ), .CI(
        \intadd_61/n4 ), .CO(\intadd_61/n3 ), .S(\intadd_51/A[2] ) );
  FA_X1 \intadd_61/U3  ( .A(\intadd_61/A[2] ), .B(\intadd_61/B[2] ), .CI(
        \intadd_61/n3 ), .CO(\intadd_61/n2 ), .S(\intadd_51/A[3] ) );
  FA_X1 \intadd_61/U2  ( .A(\intadd_61/A[3] ), .B(\intadd_61/B[3] ), .CI(
        \intadd_61/n2 ), .CO(\intadd_61/n1 ), .S(\intadd_51/A[4] ) );
  FA_X1 \intadd_62/U5  ( .A(\intadd_62/A[0] ), .B(\intadd_62/B[0] ), .CI(n2196), .CO(\intadd_62/n4 ), .S(\intadd_52/A[1] ) );
  FA_X1 \intadd_62/U4  ( .A(\intadd_62/A[1] ), .B(\intadd_62/B[1] ), .CI(
        \intadd_62/n4 ), .CO(\intadd_62/n3 ), .S(\intadd_52/B[2] ) );
  FA_X1 \intadd_62/U3  ( .A(\intadd_62/A[2] ), .B(\intadd_62/B[2] ), .CI(
        \intadd_62/n3 ), .CO(\intadd_62/n2 ), .S(\intadd_52/B[3] ) );
  FA_X1 \intadd_62/U2  ( .A(\intadd_62/A[3] ), .B(\intadd_62/B[3] ), .CI(
        \intadd_62/n2 ), .CO(\intadd_62/n1 ), .S(\intadd_52/B[4] ) );
  FA_X1 \intadd_63/U5  ( .A(\intadd_63/A[0] ), .B(\intadd_63/B[0] ), .CI(
        \intadd_63/CI ), .CO(\intadd_63/n4 ), .S(\intadd_63/SUM[0] ) );
  FA_X1 \intadd_63/U4  ( .A(\intadd_63/A[1] ), .B(\intadd_63/B[1] ), .CI(
        \intadd_63/n4 ), .CO(\intadd_63/n3 ), .S(\intadd_63/SUM[1] ) );
  FA_X1 \intadd_63/U3  ( .A(\intadd_49/SUM[0] ), .B(\intadd_63/B[2] ), .CI(
        \intadd_63/n3 ), .CO(\intadd_63/n2 ), .S(\intadd_61/A[3] ) );
  FA_X1 \intadd_63/U2  ( .A(\intadd_50/SUM[2] ), .B(\intadd_63/B[3] ), .CI(
        \intadd_63/n2 ), .CO(\intadd_63/n1 ), .S(\intadd_63/SUM[3] ) );
  FA_X1 \intadd_64/U5  ( .A(\intadd_64/A[0] ), .B(\intadd_64/B[0] ), .CI(
        \intadd_64/CI ), .CO(\intadd_64/n4 ), .S(\intadd_46/B[1] ) );
  FA_X1 \intadd_64/U4  ( .A(\intadd_64/A[1] ), .B(\intadd_64/B[1] ), .CI(
        \intadd_64/n4 ), .CO(\intadd_64/n3 ), .S(\intadd_46/B[2] ) );
  FA_X1 \intadd_64/U3  ( .A(\intadd_64/A[2] ), .B(\intadd_64/B[2] ), .CI(
        \intadd_64/n3 ), .CO(\intadd_64/n2 ), .S(\intadd_64/SUM[2] ) );
  FA_X1 \intadd_64/U2  ( .A(\intadd_64/A[3] ), .B(\intadd_64/B[3] ), .CI(
        \intadd_64/n2 ), .CO(\intadd_64/n1 ), .S(\intadd_46/A[4] ) );
  FA_X1 \intadd_65/U5  ( .A(\intadd_65/A[0] ), .B(\intadd_65/B[0] ), .CI(
        \intadd_65/CI ), .CO(\intadd_65/n4 ), .S(\intadd_65/SUM[0] ) );
  FA_X1 \intadd_65/U4  ( .A(\intadd_65/A[1] ), .B(\intadd_65/B[1] ), .CI(
        \intadd_65/n4 ), .CO(\intadd_65/n3 ), .S(\intadd_65/SUM[1] ) );
  FA_X1 \intadd_65/U3  ( .A(\intadd_65/A[2] ), .B(\intadd_65/B[2] ), .CI(
        \intadd_65/n3 ), .CO(\intadd_65/n2 ), .S(\intadd_65/SUM[2] ) );
  FA_X1 \intadd_65/U2  ( .A(\intadd_65/A[3] ), .B(\intadd_65/B[3] ), .CI(
        \intadd_65/n2 ), .CO(\intadd_65/n1 ), .S(\intadd_65/SUM[3] ) );
  FA_X1 \intadd_66/U5  ( .A(\intadd_66/A[0] ), .B(\intadd_66/B[0] ), .CI(
        \intadd_66/CI ), .CO(\intadd_66/n4 ), .S(\intadd_64/B[2] ) );
  FA_X1 \intadd_66/U4  ( .A(\intadd_66/A[1] ), .B(\intadd_66/B[1] ), .CI(
        \intadd_66/n4 ), .CO(\intadd_66/n3 ), .S(\intadd_64/A[3] ) );
  FA_X1 \intadd_66/U3  ( .A(\intadd_66/A[2] ), .B(\intadd_66/B[2] ), .CI(
        \intadd_66/n3 ), .CO(\intadd_66/n2 ), .S(\intadd_66/SUM[2] ) );
  FA_X1 \intadd_66/U2  ( .A(\intadd_66/A[3] ), .B(\intadd_65/SUM[2] ), .CI(
        \intadd_66/n2 ), .CO(\intadd_66/n1 ), .S(\intadd_66/SUM[3] ) );
  FA_X1 \intadd_67/U5  ( .A(\intadd_67/A[0] ), .B(\intadd_67/B[0] ), .CI(
        \intadd_67/CI ), .CO(\intadd_67/n4 ), .S(\intadd_67/SUM[0] ) );
  FA_X1 \intadd_67/U4  ( .A(\intadd_67/A[1] ), .B(\intadd_67/B[1] ), .CI(
        \intadd_67/n4 ), .CO(\intadd_67/n3 ), .S(\intadd_67/SUM[1] ) );
  FA_X1 \intadd_67/U3  ( .A(\intadd_67/A[2] ), .B(\intadd_67/B[2] ), .CI(
        \intadd_67/n3 ), .CO(\intadd_67/n2 ), .S(\intadd_67/SUM[2] ) );
  FA_X1 \intadd_67/U2  ( .A(\intadd_67/A[3] ), .B(\intadd_56/SUM[1] ), .CI(
        \intadd_67/n2 ), .CO(\intadd_67/n1 ), .S(\intadd_67/SUM[3] ) );
  FA_X1 \intadd_68/U5  ( .A(\intadd_68/A[0] ), .B(n2187), .CI(\intadd_68/CI ), 
        .CO(\intadd_68/n4 ), .S(\intadd_68/SUM[0] ) );
  FA_X1 \intadd_68/U4  ( .A(\intadd_68/A[1] ), .B(\intadd_68/B[1] ), .CI(
        \intadd_68/n4 ), .CO(\intadd_68/n3 ), .S(\intadd_68/SUM[1] ) );
  FA_X1 \intadd_68/U3  ( .A(\intadd_68/A[2] ), .B(\intadd_68/B[2] ), .CI(
        \intadd_68/n3 ), .CO(\intadd_68/n2 ), .S(\intadd_68/SUM[2] ) );
  FA_X1 \intadd_68/U2  ( .A(\intadd_68/A[3] ), .B(\intadd_68/B[3] ), .CI(
        \intadd_68/n2 ), .CO(\intadd_68/n1 ), .S(\intadd_68/SUM[3] ) );
  FA_X1 \intadd_69/U5  ( .A(\intadd_69/A[0] ), .B(n2188), .CI(\intadd_69/CI ), 
        .CO(\intadd_69/n4 ), .S(\intadd_69/SUM[0] ) );
  FA_X1 \intadd_69/U4  ( .A(\intadd_69/A[1] ), .B(\intadd_69/B[1] ), .CI(
        \intadd_69/n4 ), .CO(\intadd_69/n3 ), .S(\intadd_69/SUM[1] ) );
  FA_X1 \intadd_69/U3  ( .A(\intadd_69/A[2] ), .B(\intadd_69/B[2] ), .CI(
        \intadd_69/n3 ), .CO(\intadd_69/n2 ), .S(\intadd_69/SUM[2] ) );
  FA_X1 \intadd_69/U2  ( .A(\intadd_69/A[3] ), .B(\intadd_68/SUM[2] ), .CI(
        \intadd_69/n2 ), .CO(\intadd_69/n1 ), .S(\intadd_69/SUM[3] ) );
  FA_X1 \intadd_70/U4  ( .A(\intadd_70/A[0] ), .B(\intadd_70/B[0] ), .CI(
        \intadd_70/CI ), .CO(\intadd_70/n3 ), .S(\intadd_53/B[1] ) );
  FA_X1 \intadd_70/U3  ( .A(\intadd_70/A[1] ), .B(\intadd_70/B[1] ), .CI(
        \intadd_70/n3 ), .CO(\intadd_70/n2 ), .S(\intadd_53/B[2] ) );
  FA_X1 \intadd_70/U2  ( .A(\intadd_70/A[2] ), .B(\intadd_70/B[2] ), .CI(
        \intadd_70/n2 ), .CO(\intadd_70/n1 ), .S(\intadd_53/B[3] ) );
  FA_X1 \intadd_71/U4  ( .A(\intadd_71/A[0] ), .B(n2183), .CI(\intadd_71/CI ), 
        .CO(\intadd_71/n3 ), .S(\intadd_71/SUM[0] ) );
  FA_X1 \intadd_71/U3  ( .A(\intadd_71/A[1] ), .B(\intadd_71/B[1] ), .CI(
        \intadd_71/n3 ), .CO(\intadd_71/n2 ), .S(\intadd_71/SUM[1] ) );
  FA_X1 \intadd_71/U2  ( .A(\intadd_47/SUM[1] ), .B(\intadd_71/B[2] ), .CI(
        \intadd_71/n2 ), .CO(\intadd_71/n1 ), .S(\intadd_71/SUM[2] ) );
  FA_X1 \intadd_72/U4  ( .A(\intadd_72/A[0] ), .B(\intadd_72/B[0] ), .CI(
        \intadd_72/CI ), .CO(\intadd_72/n3 ), .S(\intadd_72/SUM[0] ) );
  FA_X1 \intadd_72/U2  ( .A(\intadd_72/A[2] ), .B(\intadd_72/B[2] ), .CI(
        \intadd_72/n2 ), .CO(\intadd_72/n1 ), .S(\intadd_72/SUM[2] ) );
  FA_X1 \intadd_73/U4  ( .A(\intadd_73/A[0] ), .B(\intadd_73/B[0] ), .CI(
        \intadd_73/CI ), .CO(\intadd_73/n3 ), .S(\intadd_73/SUM[0] ) );
  FA_X1 \intadd_73/U3  ( .A(\intadd_73/A[1] ), .B(\intadd_73/B[1] ), .CI(
        \intadd_73/n3 ), .CO(\intadd_73/n2 ), .S(\intadd_73/SUM[1] ) );
  FA_X1 \intadd_73/U2  ( .A(\intadd_51/SUM[1] ), .B(\intadd_73/B[2] ), .CI(
        \intadd_73/n2 ), .CO(\intadd_73/n1 ), .S(\intadd_62/A[3] ) );
  FA_X1 \intadd_74/U4  ( .A(\intadd_74/A[0] ), .B(\intadd_74/B[0] ), .CI(
        \intadd_74/CI ), .CO(\intadd_74/n3 ), .S(\intadd_74/SUM[0] ) );
  FA_X1 \intadd_74/U3  ( .A(\intadd_74/A[1] ), .B(\intadd_74/B[1] ), .CI(
        \intadd_74/n3 ), .CO(\intadd_74/n2 ), .S(\intadd_74/SUM[1] ) );
  FA_X1 \intadd_74/U2  ( .A(\intadd_74/A[2] ), .B(\intadd_74/B[2] ), .CI(
        \intadd_74/n2 ), .CO(\intadd_74/n1 ), .S(\intadd_74/SUM[2] ) );
  FA_X1 \intadd_75/U4  ( .A(\intadd_75/A[0] ), .B(\intadd_75/B[0] ), .CI(
        \intadd_75/CI ), .CO(\intadd_75/n3 ), .S(\intadd_75/SUM[0] ) );
  FA_X1 \intadd_75/U3  ( .A(\intadd_75/A[1] ), .B(\intadd_75/B[1] ), .CI(
        \intadd_75/n3 ), .CO(\intadd_75/n2 ), .S(\intadd_75/SUM[1] ) );
  FA_X1 \intadd_75/U2  ( .A(\intadd_75/A[2] ), .B(\intadd_65/SUM[0] ), .CI(
        \intadd_75/n2 ), .CO(\intadd_75/n1 ), .S(\intadd_64/B[3] ) );
  FA_X1 \intadd_76/U4  ( .A(\intadd_76/A[0] ), .B(\intadd_76/B[0] ), .CI(
        \intadd_76/CI ), .CO(\intadd_76/n3 ), .S(\intadd_76/SUM[0] ) );
  FA_X1 \intadd_76/U3  ( .A(\intadd_76/A[1] ), .B(\intadd_76/B[1] ), .CI(
        \intadd_76/n3 ), .CO(\intadd_76/n2 ), .S(\intadd_76/SUM[1] ) );
  FA_X1 \intadd_76/U2  ( .A(\intadd_76/A[2] ), .B(\intadd_76/B[2] ), .CI(
        \intadd_76/n2 ), .CO(\intadd_76/n1 ), .S(\intadd_76/SUM[2] ) );
  FA_X1 \intadd_77/U4  ( .A(\intadd_77/A[0] ), .B(\intadd_77/B[0] ), .CI(
        \intadd_55/SUM[0] ), .CO(\intadd_77/n3 ), .S(\intadd_65/A[3] ) );
  FA_X1 \intadd_77/U3  ( .A(\intadd_77/A[1] ), .B(\intadd_55/SUM[1] ), .CI(
        \intadd_77/n3 ), .CO(\intadd_77/n2 ), .S(\intadd_77/SUM[1] ) );
  FA_X1 \intadd_77/U2  ( .A(\intadd_67/SUM[3] ), .B(\intadd_55/SUM[2] ), .CI(
        \intadd_77/n2 ), .CO(\intadd_77/n1 ), .S(\intadd_77/SUM[2] ) );
  FA_X1 \intadd_78/U4  ( .A(\intadd_78/A[0] ), .B(\intadd_78/B[0] ), .CI(
        \intadd_78/CI ), .CO(\intadd_78/n3 ), .S(\intadd_78/SUM[0] ) );
  FA_X1 \intadd_78/U3  ( .A(\intadd_78/A[1] ), .B(\intadd_78/B[1] ), .CI(
        \intadd_78/n3 ), .CO(\intadd_78/n2 ), .S(\intadd_78/SUM[1] ) );
  FA_X1 \intadd_78/U2  ( .A(\intadd_78/A[2] ), .B(\intadd_78/B[2] ), .CI(
        \intadd_78/n2 ), .CO(\intadd_78/n1 ), .S(\intadd_78/SUM[2] ) );
  FA_X1 \intadd_79/U4  ( .A(\intadd_79/A[0] ), .B(\intadd_79/B[0] ), .CI(
        \intadd_79/CI ), .CO(\intadd_79/n3 ), .S(\intadd_79/SUM[0] ) );
  FA_X1 \intadd_79/U3  ( .A(\intadd_53/SUM[0] ), .B(\intadd_79/B[1] ), .CI(
        \intadd_79/n3 ), .CO(\intadd_79/n2 ), .S(\intadd_56/B[3] ) );
  FA_X1 \intadd_79/U2  ( .A(\intadd_79/A[2] ), .B(\intadd_79/B[2] ), .CI(
        \intadd_79/n2 ), .CO(\intadd_79/n1 ), .S(\intadd_56/B[4] ) );
  FA_X1 \intadd_80/U4  ( .A(\intadd_80/A[0] ), .B(\intadd_80/B[0] ), .CI(
        \intadd_80/CI ), .CO(\intadd_80/n3 ), .S(\intadd_78/A[0] ) );
  FA_X1 \intadd_80/U3  ( .A(\intadd_80/A[1] ), .B(\intadd_80/B[1] ), .CI(
        \intadd_80/n3 ), .CO(\intadd_80/n2 ), .S(\intadd_78/B[1] ) );
  FA_X1 \intadd_80/U2  ( .A(\intadd_80/A[2] ), .B(\intadd_80/B[2] ), .CI(
        \intadd_80/n2 ), .CO(\intadd_80/n1 ), .S(\intadd_78/A[2] ) );
  FA_X1 \intadd_81/U4  ( .A(\intadd_81/A[0] ), .B(\intadd_81/B[0] ), .CI(
        \intadd_81/CI ), .CO(\intadd_81/n3 ), .S(\intadd_81/SUM[0] ) );
  FA_X1 \intadd_81/U3  ( .A(\intadd_69/SUM[0] ), .B(\intadd_81/B[1] ), .CI(
        \intadd_81/n3 ), .CO(\intadd_81/n2 ), .S(\intadd_60/B[3] ) );
  FA_X1 \intadd_81/U2  ( .A(\intadd_68/SUM[0] ), .B(\intadd_81/B[2] ), .CI(
        \intadd_81/n2 ), .CO(\intadd_81/n1 ), .S(\intadd_81/SUM[2] ) );
  INV_X1 U4 ( .A(a[9]), .ZN(n1250) );
  AND2_X1 U5 ( .A1(n1706), .A2(a[13]), .ZN(\intadd_69/A[0] ) );
  INV_X1 U8 ( .A(\intadd_56/SUM[2] ), .ZN(n356) );
  INV_X1 U9 ( .A(\intadd_78/SUM[0] ), .ZN(\intadd_55/B[3] ) );
  INV_X1 U10 ( .A(\intadd_80/n1 ), .ZN(\intadd_53/A[2] ) );
  INV_X1 U13 ( .A(n2106), .ZN(n2104) );
  AND2_X1 U14 ( .A1(\intadd_50/n1 ), .A2(\intadd_49/SUM[4] ), .ZN(n2111) );
  INV_X1 U16 ( .A(a[5]), .ZN(n1180) );
  INV_X1 U19 ( .A(a[7]), .ZN(n1024) );
  INV_X1 U20 ( .A(n1712), .ZN(n1752) );
  INV_X1 U21 ( .A(n1618), .ZN(n1596) );
  AND2_X1 U25 ( .A1(n400), .A2(n401), .ZN(n1068) );
  INV_X1 U26 ( .A(b[14]), .ZN(n1602) );
  INV_X1 U27 ( .A(n1529), .ZN(n1437) );
  INV_X1 U29 ( .A(\intadd_79/SUM[0] ), .ZN(\intadd_78/B[0] ) );
  INV_X1 U30 ( .A(n482), .ZN(n483) );
  INV_X1 U31 ( .A(n649), .ZN(n181) );
  OR2_X1 U32 ( .A1(n110), .A2(n109), .ZN(n103) );
  AND2_X1 U33 ( .A1(n1691), .A2(n1690), .ZN(n1644) );
  INV_X1 U34 ( .A(n641), .ZN(\intadd_65/A[2] ) );
  OR2_X1 U36 ( .A1(n363), .A2(n362), .ZN(n364) );
  INV_X1 U38 ( .A(\intadd_74/SUM[1] ), .ZN(\intadd_46/A[2] ) );
  INV_X1 U39 ( .A(\intadd_74/n1 ), .ZN(n333) );
  AND2_X1 U40 ( .A1(n2092), .A2(n338), .ZN(n351) );
  INV_X1 U41 ( .A(\intadd_76/n1 ), .ZN(n353) );
  INV_X1 U44 ( .A(n1423), .ZN(n1424) );
  INV_X1 U45 ( .A(n580), .ZN(n382) );
  INV_X1 U47 ( .A(n1916), .ZN(n600) );
  INV_X1 U48 ( .A(n1933), .ZN(n601) );
  OR2_X1 U49 ( .A1(n2026), .A2(n1930), .ZN(n2029) );
  INV_X1 U52 ( .A(n1697), .ZN(n1738) );
  INV_X1 U53 ( .A(n1883), .ZN(n1375) );
  INV_X1 U54 ( .A(a[11]), .ZN(n124) );
  OR2_X1 U55 ( .A1(a[9]), .A2(a[10]), .ZN(n125) );
  INV_X1 U56 ( .A(a[2]), .ZN(n475) );
  INV_X1 U57 ( .A(n213), .ZN(n782) );
  INV_X1 U58 ( .A(a[17]), .ZN(n215) );
  AND2_X1 U59 ( .A1(n1183), .A2(a[5]), .ZN(\intadd_49/B[0] ) );
  INV_X1 U62 ( .A(n1852), .ZN(n1766) );
  INV_X1 U64 ( .A(n1742), .ZN(n1666) );
  AND2_X1 U65 ( .A1(n125), .A2(b[0]), .ZN(n1729) );
  INV_X1 U67 ( .A(n1481), .ZN(n1580) );
  INV_X1 U68 ( .A(n1627), .ZN(n1629) );
  AND2_X1 U70 ( .A1(n1549), .A2(n1548), .ZN(n1543) );
  AND2_X1 U71 ( .A1(n752), .A2(n751), .ZN(n766) );
  INV_X1 U76 ( .A(n1409), .ZN(n1574) );
  INV_X1 U77 ( .A(b[7]), .ZN(n1735) );
  INV_X1 U79 ( .A(a[13]), .ZN(n232) );
  INV_X1 U81 ( .A(b[4]), .ZN(n1651) );
  INV_X1 U83 ( .A(n1725), .ZN(n1703) );
  INV_X1 U85 ( .A(n1701), .ZN(n1741) );
  INV_X1 U88 ( .A(n1722), .ZN(n1689) );
  INV_X1 U91 ( .A(b[13]), .ZN(n1670) );
  INV_X1 U98 ( .A(a[19]), .ZN(n1442) );
  INV_X1 U100 ( .A(n1231), .ZN(n1289) );
  OR2_X1 U104 ( .A1(n90), .A2(n1742), .ZN(n93) );
  AND2_X1 U108 ( .A1(n648), .A2(n647), .ZN(n652) );
  INV_X1 U111 ( .A(n73), .ZN(n1760) );
  INV_X1 U112 ( .A(n1659), .ZN(n1631) );
  INV_X1 U113 ( .A(n1562), .ZN(n1568) );
  INV_X1 U115 ( .A(n1585), .ZN(n1587) );
  INV_X1 U117 ( .A(n1460), .ZN(n1500) );
  INV_X1 U119 ( .A(n1269), .ZN(n1270) );
  INV_X1 U120 ( .A(n1617), .ZN(n1276) );
  INV_X1 U121 ( .A(n1389), .ZN(n1619) );
  INV_X1 U122 ( .A(b[10]), .ZN(n1732) );
  INV_X1 U126 ( .A(\intadd_52/SUM[0] ), .ZN(\intadd_80/A[2] ) );
  INV_X1 U127 ( .A(n137), .ZN(n138) );
  INV_X1 U128 ( .A(n1215), .ZN(n1219) );
  INV_X1 U129 ( .A(\intadd_77/n1 ), .ZN(n360) );
  AND2_X1 U130 ( .A1(n1200), .A2(n1199), .ZN(n1202) );
  OR2_X1 U131 ( .A1(\intadd_71/SUM[0] ), .A2(n404), .ZN(n406) );
  INV_X1 U132 ( .A(n620), .ZN(\intadd_47/A[1] ) );
  INV_X1 U133 ( .A(b[20]), .ZN(n1309) );
  INV_X1 U134 ( .A(n1394), .ZN(n1528) );
  INV_X1 U135 ( .A(n190), .ZN(n1377) );
  INV_X1 U137 ( .A(b[21]), .ZN(n1991) );
  AND2_X1 U138 ( .A1(a[1]), .A2(a[2]), .ZN(n1330) );
  INV_X1 U139 ( .A(a[3]), .ZN(n1331) );
  OR2_X1 U141 ( .A1(n1826), .A2(n2051), .ZN(n1832) );
  INV_X1 U142 ( .A(\intadd_75/SUM[0] ), .ZN(\intadd_74/B[1] ) );
  INV_X1 U143 ( .A(\intadd_46/SUM[1] ), .ZN(n1839) );
  INV_X1 U145 ( .A(n371), .ZN(n375) );
  INV_X1 U146 ( .A(n1348), .ZN(n1351) );
  INV_X1 U147 ( .A(\intadd_73/SUM[1] ), .ZN(n1353) );
  INV_X1 U148 ( .A(n1420), .ZN(n1354) );
  OR2_X1 U149 ( .A1(n558), .A2(n557), .ZN(n561) );
  INV_X1 U150 ( .A(\intadd_63/n1 ), .ZN(n582) );
  AND2_X1 U151 ( .A1(n1917), .A2(n1915), .ZN(n592) );
  INV_X1 U155 ( .A(b[22]), .ZN(n1996) );
  INV_X1 U157 ( .A(b[18]), .ZN(n1247) );
  INV_X1 U158 ( .A(a[23]), .ZN(n2167) );
  INV_X1 U159 ( .A(n2137), .ZN(n2150) );
  OR2_X1 U160 ( .A1(n2140), .A2(n2142), .ZN(n2149) );
  INV_X1 U161 ( .A(a[1]), .ZN(n1205) );
  INV_X1 U165 ( .A(n335), .ZN(n2092) );
  OR2_X1 U166 ( .A1(\intadd_46/A[4] ), .A2(n333), .ZN(n334) );
  INV_X1 U167 ( .A(\intadd_76/SUM[0] ), .ZN(\intadd_66/A[3] ) );
  INV_X1 U169 ( .A(\intadd_65/n1 ), .ZN(n1903) );
  INV_X1 U171 ( .A(\intadd_78/SUM[1] ), .ZN(\intadd_55/B[4] ) );
  INV_X1 U172 ( .A(\intadd_78/SUM[2] ), .ZN(\intadd_56/A[4] ) );
  AND2_X1 U174 ( .A1(n2068), .A2(n2070), .ZN(n1952) );
  AND2_X1 U178 ( .A1(n2076), .A2(n2103), .ZN(n2077) );
  AND2_X1 U180 ( .A1(\intadd_48/SUM[4] ), .A2(\intadd_47/n1 ), .ZN(n1988) );
  INV_X1 U181 ( .A(n1920), .ZN(n1922) );
  INV_X1 U182 ( .A(n2146), .ZN(n2037) );
  INV_X1 U185 ( .A(n1981), .ZN(n1911) );
  INV_X1 U186 ( .A(n1946), .ZN(n1949) );
  OR2_X1 U187 ( .A1(\intadd_52/n1 ), .A2(n574), .ZN(n2071) );
  INV_X1 U188 ( .A(n1965), .ZN(n2017) );
  INV_X1 U189 ( .A(n1960), .ZN(n2078) );
  INV_X1 U190 ( .A(n2126), .ZN(n2120) );
  INV_X1 U191 ( .A(n2148), .ZN(n1938) );
  INV_X1 U192 ( .A(n2156), .ZN(n2158) );
  INV_X1 U193 ( .A(n611), .ZN(\intadd_58/B[3] ) );
  OR2_X1 U194 ( .A1(n2035), .A2(n2034), .ZN(\d[41]_BAR ) );
  XOR2_X1 U195 ( .A(n108), .B(n107), .Z(\d[6]_BAR ) );
  INV_X1 U197 ( .A(b[5]), .ZN(n1611) );
  INV_X1 U198 ( .A(n144), .ZN(n1861) );
  NOR2_X1 U199 ( .A1(\intadd_58/SUM[0] ), .A2(n322), .ZN(n2) );
  INV_X1 U200 ( .A(n1902), .ZN(n1262) );
  INV_X1 U202 ( .A(b[23]), .ZN(n2165) );
  INV_X1 U203 ( .A(n1862), .ZN(n1599) );
  INV_X1 U204 ( .A(b[11]), .ZN(n1717) );
  XOR2_X1 U205 ( .A(\intadd_54/n3 ), .B(n111), .Z(\d[11]_BAR ) );
  INV_X1 U206 ( .A(n1999), .ZN(n1287) );
  INV_X1 U207 ( .A(n450), .ZN(n448) );
  INV_X1 U209 ( .A(n1308), .ZN(n1206) );
  INV_X1 U210 ( .A(n1171), .ZN(n1173) );
  INV_X1 U212 ( .A(n1119), .ZN(n1115) );
  INV_X1 U213 ( .A(n615), .ZN(n616) );
  INV_X1 U214 ( .A(n400), .ZN(n403) );
  INV_X1 U215 ( .A(b[9]), .ZN(n1684) );
  INV_X1 U216 ( .A(b[19]), .ZN(n1341) );
  INV_X1 U217 ( .A(n1804), .ZN(n87) );
  INV_X1 U218 ( .A(n1856), .ZN(n1865) );
  INV_X1 U219 ( .A(n1745), .ZN(n1709) );
  INV_X1 U220 ( .A(n1718), .ZN(n1681) );
  INV_X1 U221 ( .A(n1707), .ZN(n650) );
  INV_X1 U222 ( .A(n1637), .ZN(n788) );
  INV_X1 U223 ( .A(n1251), .ZN(n63) );
  INV_X1 U225 ( .A(n1439), .ZN(n1450) );
  INV_X1 U226 ( .A(n1531), .ZN(n1435) );
  INV_X1 U227 ( .A(n1368), .ZN(n1336) );
  INV_X1 U228 ( .A(n1300), .ZN(n1361) );
  INV_X1 U232 ( .A(b[12]), .ZN(n1273) );
  INV_X1 U233 ( .A(n1108), .ZN(n1106) );
  INV_X1 U234 ( .A(n1174), .ZN(n1146) );
  INV_X1 U235 ( .A(n1137), .ZN(n1141) );
  INV_X1 U236 ( .A(n1769), .ZN(n1753) );
  INV_X1 U238 ( .A(n953), .ZN(n897) );
  INV_X1 U239 ( .A(n925), .ZN(n905) );
  INV_X1 U240 ( .A(n833), .ZN(n1579) );
  INV_X1 U241 ( .A(n914), .ZN(n225) );
  INV_X1 U242 ( .A(b[15]), .ZN(n1131) );
  INV_X1 U243 ( .A(n848), .ZN(n835) );
  INV_X1 U244 ( .A(a[15]), .ZN(n633) );
  INV_X1 U245 ( .A(n1183), .ZN(n17) );
  INV_X1 U246 ( .A(n1847), .ZN(n96) );
  INV_X1 U248 ( .A(n1672), .ZN(n639) );
  INV_X1 U250 ( .A(n1633), .ZN(n779) );
  INV_X1 U252 ( .A(n776), .ZN(n1510) );
  INV_X1 U253 ( .A(b[6]), .ZN(n1859) );
  INV_X1 U255 ( .A(n1370), .ZN(n1339) );
  INV_X1 U256 ( .A(n1316), .ZN(n1293) );
  INV_X1 U257 ( .A(n1770), .ZN(n1715) );
  INV_X1 U258 ( .A(b[8]), .ZN(n1694) );
  INV_X1 U259 ( .A(n1167), .ZN(n1169) );
  INV_X1 U261 ( .A(n1080), .ZN(n1084) );
  INV_X1 U262 ( .A(n1123), .ZN(n404) );
  INV_X1 U263 ( .A(n1022), .ZN(n991) );
  INV_X1 U264 ( .A(n943), .ZN(n936) );
  INV_X1 U265 ( .A(n927), .ZN(n907) );
  INV_X1 U266 ( .A(n251), .ZN(n252) );
  INV_X1 U267 ( .A(n808), .ZN(n296) );
  INV_X1 U269 ( .A(n2000), .ZN(n2001) );
  INV_X1 U270 ( .A(n1632), .ZN(n780) );
  INV_X1 U271 ( .A(n1586), .ZN(n1584) );
  INV_X1 U273 ( .A(n1592), .ZN(n1515) );
  INV_X1 U274 ( .A(b[3]), .ZN(n1787) );
  INV_X1 U276 ( .A(n1356), .ZN(n1357) );
  INV_X1 U277 ( .A(n1216), .ZN(n1218) );
  INV_X1 U278 ( .A(n1319), .ZN(n1277) );
  INV_X1 U279 ( .A(\intadd_63/SUM[1] ), .ZN(n1163) );
  INV_X1 U280 ( .A(\intadd_49/SUM[1] ), .ZN(n1100) );
  INV_X1 U281 ( .A(n921), .ZN(n902) );
  INV_X1 U282 ( .A(n844), .ZN(n827) );
  INV_X1 U285 ( .A(b[2]), .ZN(n1740) );
  INV_X1 U287 ( .A(\intadd_72/SUM[0] ), .ZN(n37) );
  INV_X1 U288 ( .A(n1828), .ZN(n1831) );
  INV_X1 U289 ( .A(n2053), .ZN(n1833) );
  INV_X1 U290 ( .A(n346), .ZN(n347) );
  INV_X1 U291 ( .A(n1575), .ZN(n1410) );
  INV_X1 U292 ( .A(n1493), .ZN(n1487) );
  INV_X1 U293 ( .A(n1498), .ZN(n1463) );
  INV_X1 U294 ( .A(n588), .ZN(n374) );
  INV_X1 U296 ( .A(n1919), .ZN(n593) );
  INV_X1 U297 ( .A(n2145), .ZN(n2147) );
  INV_X1 U298 ( .A(n1449), .ZN(n1900) );
  INV_X1 U300 ( .A(a[21]), .ZN(n130) );
  INV_X1 U301 ( .A(n1327), .ZN(n1176) );
  INV_X1 U302 ( .A(n369), .ZN(n177) );
  INV_X1 U303 ( .A(n1496), .ZN(n1468) );
  INV_X1 U304 ( .A(n2062), .ZN(n373) );
  INV_X1 U305 ( .A(n2103), .ZN(n1956) );
  INV_X1 U306 ( .A(\intadd_68/SUM[1] ), .ZN(n207) );
  INV_X1 U308 ( .A(n1924), .ZN(n604) );
  INV_X1 U309 ( .A(n2161), .ZN(n2006) );
  INV_X1 U311 ( .A(n2051), .ZN(n1977) );
  INV_X1 U313 ( .A(\intadd_60/SUM[3] ), .ZN(n2118) );
  INV_X1 U314 ( .A(n1992), .ZN(n1886) );
  INV_X1 U316 ( .A(n8), .ZN(n9) );
  INV_X1 U317 ( .A(n25), .ZN(n2043) );
  INV_X1 U318 ( .A(n2122), .ZN(n2123) );
  INV_X1 U319 ( .A(n1950), .ZN(n1929) );
  INV_X1 U321 ( .A(b[1]), .ZN(n2086) );
  INV_X1 U322 ( .A(n1908), .ZN(n1909) );
  NAND2_X1 U324 ( .A1(a[4]), .A2(a[3]), .ZN(n1183) );
  NOR2_X1 U325 ( .A1(a[2]), .A2(a[1]), .ZN(n1327) );
  NOR2_X1 U326 ( .A1(n1330), .A2(n1327), .ZN(n8) );
  MUX2_X1 U327 ( .A(n1850), .B(n1849), .S(b[1]), .Z(n5) );
  NAND2_X1 U328 ( .A1(n1327), .A2(a[3]), .ZN(n1852) );
  NOR2_X1 U329 ( .A1(n475), .A2(a[3]), .ZN(n1171) );
  MUX2_X1 U330 ( .A(n1852), .B(n1851), .S(b[0]), .Z(n4) );
  NAND2_X1 U331 ( .A1(n5), .A2(n4), .ZN(n24) );
  NAND2_X1 U332 ( .A1(a[1]), .A2(a[0]), .ZN(n1856) );
  NAND2_X1 U336 ( .A1(n24), .A2(n23), .ZN(n25) );
  AOI21_X1 U337 ( .B1(a[1]), .B2(n2086), .A(n1867), .ZN(n2085) );
  MUX2_X1 U338 ( .A(n2085), .B(n9), .S(b[0]), .Z(n1936) );
  MUX2_X1 U339 ( .A(n1856), .B(n1855), .S(b[2]), .Z(n11) );
  NAND2_X1 U340 ( .A1(n1867), .A2(n2086), .ZN(n10) );
  AND2_X1 U341 ( .A1(n11), .A2(n10), .ZN(n1935) );
  NOR2_X1 U342 ( .A1(n1936), .A2(n1935), .ZN(n22) );
  OR2_X1 U344 ( .A1(n1330), .A2(b[0]), .ZN(n12) );
  AOI21_X1 U345 ( .B1(n12), .B2(n1176), .A(n1331), .ZN(n21) );
  NAND2_X1 U347 ( .A1(n2043), .A2(n2047), .ZN(n1970) );
  INV_X1 U348 ( .A(n1970), .ZN(n33) );
  NAND2_X1 U352 ( .A1(n38), .A2(b[0]), .ZN(n42) );
  NOR2_X1 U353 ( .A1(n42), .A2(n17), .ZN(n28) );
  XOR2_X1 U354 ( .A(n27), .B(n28), .Z(n20) );
  MUX2_X1 U355 ( .A(n1850), .B(n1849), .S(b[2]), .Z(n19) );
  MUX2_X1 U356 ( .A(n1852), .B(n1851), .S(b[1]), .Z(n18) );
  NAND2_X1 U357 ( .A1(n19), .A2(n18), .ZN(n26) );
  XOR2_X1 U358 ( .A(n20), .B(n26), .Z(n2044) );
  NOR2_X1 U359 ( .A1(n22), .A2(n21), .ZN(n2045) );
  NOR2_X1 U360 ( .A1(n24), .A2(n23), .ZN(n1968) );
  OAI21_X1 U361 ( .B1(n2045), .B2(n1968), .A(n25), .ZN(n34) );
  NAND2_X1 U363 ( .A1(n27), .A2(n28), .ZN(n31) );
  OAI211_X1 U367 ( .C1(n33), .C2(n2044), .A(n34), .B(n1972), .ZN(n36) );
  NAND2_X1 U368 ( .A1(n2044), .A2(n34), .ZN(n1971) );
  AOI22_X1 U369 ( .A1(n37), .A2(n36), .B1(n1971), .B2(n35), .ZN(n107) );
  NAND3_X1 U370 ( .A1(n38), .A2(n1180), .A3(n1183), .ZN(n144) );
  MUX2_X1 U371 ( .A(n144), .B(n1788), .S(n2086), .Z(n41) );
  NOR2_X1 U372 ( .A1(n1183), .A2(a[5]), .ZN(n1862) );
  MUX2_X1 U373 ( .A(n1789), .B(n1599), .S(b[0]), .Z(n40) );
  NAND2_X1 U374 ( .A1(n41), .A2(n40), .ZN(n642) );
  AND2_X1 U375 ( .A1(n42), .A2(\intadd_49/B[0] ), .ZN(n643) );
  NAND2_X1 U376 ( .A1(n642), .A2(n643), .ZN(n1799) );
  MUX2_X1 U377 ( .A(n1850), .B(n1849), .S(b[4]), .Z(n44) );
  MUX2_X1 U378 ( .A(n1852), .B(n1851), .S(b[3]), .Z(n43) );
  NAND2_X1 U379 ( .A1(n44), .A2(n43), .ZN(n1796) );
  XOR2_X1 U380 ( .A(n1799), .B(n1796), .Z(n50) );
  XOR2_X1 U384 ( .A(a[5]), .B(a[6]), .Z(n776) );
  AND2_X1 U385 ( .A1(n776), .A2(b[0]), .ZN(n1779) );
  XNOR2_X1 U386 ( .A(n1778), .B(n1779), .ZN(n49) );
  MUX2_X1 U387 ( .A(n144), .B(n1788), .S(n1740), .Z(n48) );
  MUX2_X1 U388 ( .A(n1789), .B(n1599), .S(b[1]), .Z(n47) );
  NAND2_X1 U389 ( .A1(n48), .A2(n47), .ZN(n1780) );
  XOR2_X1 U390 ( .A(n49), .B(n1780), .Z(n1797) );
  XOR2_X1 U391 ( .A(n50), .B(n1797), .Z(n106) );
  OAI21_X1 U392 ( .B1(n107), .B2(n106), .A(\intadd_72/n3 ), .ZN(n52) );
  NAND2_X1 U393 ( .A1(n107), .A2(n106), .ZN(n51) );
  NAND2_X1 U394 ( .A1(n52), .A2(n51), .ZN(\intadd_72/n2 ) );
  MUX2_X1 U395 ( .A(n1850), .B(n1849), .S(b[7]), .Z(n54) );
  MUX2_X1 U396 ( .A(n1852), .B(n1851), .S(b[6]), .Z(n53) );
  MUX2_X1 U397 ( .A(n144), .B(n1788), .S(n1611), .Z(n56) );
  MUX2_X1 U398 ( .A(n1789), .B(n1599), .S(b[4]), .Z(n55) );
  NOR2_X1 U399 ( .A1(n1835), .A2(n60), .ZN(n62) );
  NAND2_X1 U400 ( .A1(n776), .A2(n1024), .ZN(n1770) );
  NAND2_X1 U401 ( .A1(n776), .A2(a[7]), .ZN(n1769) );
  NOR2_X1 U402 ( .A1(n1769), .A2(b[3]), .ZN(n57) );
  AOI21_X1 U403 ( .B1(b[3]), .B2(n1715), .A(n57), .ZN(n59) );
  NOR3_X1 U404 ( .A1(n1024), .A2(a[5]), .A3(a[6]), .ZN(n1712) );
  NAND2_X1 U405 ( .A1(a[6]), .A2(a[5]), .ZN(n645) );
  MUX2_X1 U406 ( .A(n1752), .B(n1751), .S(b[2]), .Z(n58) );
  NAND2_X1 U407 ( .A1(n59), .A2(n58), .ZN(n1834) );
  OAI22_X1 U409 ( .A1(n62), .A2(n1834), .B1(n1836), .B2(n61), .ZN(n81) );
  NAND2_X1 U410 ( .A1(a[8]), .A2(a[7]), .ZN(n1251) );
  NOR2_X1 U411 ( .A1(a[7]), .A2(a[8]), .ZN(n1255) );
  NOR2_X1 U412 ( .A1(n63), .A2(n1255), .ZN(n1557) );
  NAND2_X1 U413 ( .A1(n1557), .A2(n1250), .ZN(n1697) );
  MUX2_X1 U414 ( .A(n1698), .B(n1697), .S(b[2]), .Z(n65) );
  NAND2_X1 U415 ( .A1(n1255), .A2(a[9]), .ZN(n1701) );
  NOR2_X1 U416 ( .A1(n1251), .A2(a[9]), .ZN(n1742) );
  MUX2_X1 U417 ( .A(n1701), .B(n1666), .S(b[1]), .Z(n64) );
  NAND2_X1 U418 ( .A1(n65), .A2(n64), .ZN(n1759) );
  NAND2_X1 U419 ( .A1(a[9]), .A2(a[10]), .ZN(n123) );
  NAND2_X1 U420 ( .A1(n1729), .A2(n123), .ZN(n1758) );
  XOR2_X1 U421 ( .A(n1759), .B(n1758), .Z(n74) );
  INV_X1 U422 ( .A(n74), .ZN(n72) );
  NOR2_X1 U423 ( .A1(n1770), .A2(n1651), .ZN(n68) );
  NOR2_X1 U424 ( .A1(n1769), .A2(b[4]), .ZN(n67) );
  MUX2_X1 U425 ( .A(n1712), .B(n1711), .S(b[3]), .Z(n66) );
  NOR3_X1 U426 ( .A1(n68), .A2(n67), .A3(n66), .ZN(n73) );
  INV_X1 U427 ( .A(n1759), .ZN(n69) );
  NOR2_X1 U428 ( .A1(n69), .A2(n73), .ZN(n1762) );
  OAI21_X1 U429 ( .B1(n1698), .B2(b[1]), .A(n1701), .ZN(n90) );
  NOR2_X1 U431 ( .A1(n1762), .A2(n70), .ZN(n71) );
  OAI21_X1 U432 ( .B1(n72), .B2(n1760), .A(n71), .ZN(n78) );
  AOI21_X1 U435 ( .B1(n81), .B2(n78), .A(n80), .ZN(n1838) );
  XNOR2_X1 U436 ( .A(\intadd_74/SUM[0] ), .B(n1838), .ZN(n77) );
  XOR2_X1 U437 ( .A(\intadd_46/SUM[1] ), .B(n77), .Z(n110) );
  INV_X1 U438 ( .A(n78), .ZN(n79) );
  NOR2_X1 U439 ( .A1(n80), .A2(n79), .ZN(n82) );
  XNOR2_X1 U440 ( .A(n82), .B(n81), .ZN(n1843) );
  MUX2_X1 U441 ( .A(n1769), .B(n1770), .S(b[2]), .Z(n84) );
  MUX2_X1 U442 ( .A(n1752), .B(n1751), .S(b[1]), .Z(n83) );
  NAND2_X1 U443 ( .A1(n84), .A2(n83), .ZN(n1805) );
  MUX2_X1 U444 ( .A(n144), .B(n1788), .S(n1651), .Z(n86) );
  MUX2_X1 U445 ( .A(n1789), .B(n1599), .S(b[3]), .Z(n85) );
  NAND2_X1 U446 ( .A1(n86), .A2(n85), .ZN(n1806) );
  NAND2_X1 U447 ( .A1(n1557), .A2(b[0]), .ZN(n1804) );
  NAND2_X1 U450 ( .A1(n1557), .A2(n2084), .ZN(n91) );
  NAND2_X1 U451 ( .A1(n1697), .A2(n91), .ZN(n92) );
  AOI22_X1 U452 ( .A1(n93), .A2(b[0]), .B1(b[1]), .B2(n92), .ZN(n1846) );
  NAND2_X1 U453 ( .A1(n1847), .A2(n1846), .ZN(n98) );
  INV_X1 U457 ( .A(n1846), .ZN(n97) );
  AOI22_X1 U458 ( .A1(n98), .A2(n1845), .B1(n97), .B2(n96), .ZN(n1842) );
  NAND2_X1 U459 ( .A1(\intadd_46/SUM[0] ), .A2(n1842), .ZN(n101) );
  AOI22_X1 U463 ( .A1(\intadd_54/n3 ), .A2(n103), .B1(n110), .B2(n109), .ZN(
        n104) );
  INV_X2 U464 ( .A(n104), .ZN(\intadd_54/n2 ) );
  XNOR2_X1 U465 ( .A(\intadd_46/A[4] ), .B(n333), .ZN(n105) );
  XNOR2_X1 U466 ( .A(\intadd_46/n2 ), .B(n105), .ZN(\d[14]_BAR ) );
  XNOR2_X1 U467 ( .A(n106), .B(\intadd_72/n3 ), .ZN(n108) );
  XNOR2_X1 U468 ( .A(n110), .B(n109), .ZN(n111) );
  INV_X2 U469 ( .A(\intadd_57/SUM[0] ), .ZN(\d[20] ) );
  INV_X2 U470 ( .A(\intadd_57/SUM[1] ), .ZN(\d[21] ) );
  XNOR2_X1 U472 ( .A(\intadd_55/SUM[3] ), .B(\intadd_67/n1 ), .ZN(n113) );
  NAND2_X1 U473 ( .A1(n114), .A2(\intadd_56/SUM[2] ), .ZN(n359) );
  NOR2_X1 U474 ( .A1(\intadd_55/SUM[3] ), .A2(\intadd_67/n1 ), .ZN(n357) );
  NAND2_X1 U475 ( .A1(n357), .A2(\intadd_56/SUM[2] ), .ZN(n112) );
  OAI211_X1 U476 ( .C1(\intadd_56/SUM[2] ), .C2(n113), .A(n359), .B(n112), 
        .ZN(\intadd_57/B[0] ) );
  INV_X2 U478 ( .A(\intadd_78/n1 ), .ZN(n116) );
  NAND2_X1 U479 ( .A1(n116), .A2(\intadd_53/SUM[2] ), .ZN(n371) );
  NOR2_X1 U480 ( .A1(n116), .A2(\intadd_53/SUM[2] ), .ZN(n1942) );
  NOR2_X1 U481 ( .A1(n375), .A2(n1942), .ZN(n180) );
  NOR2_X1 U483 ( .A1(a[17]), .A2(a[18]), .ZN(n1453) );
  NOR2_X1 U484 ( .A1(n1443), .A2(n1453), .ZN(n1517) );
  NAND2_X1 U485 ( .A1(n215), .A2(a[19]), .ZN(n1899) );
  NOR2_X1 U486 ( .A1(n1899), .A2(a[18]), .ZN(n1439) );
  NAND2_X1 U487 ( .A1(n1439), .A2(n1651), .ZN(n119) );
  NOR2_X1 U488 ( .A1(n117), .A2(a[19]), .ZN(n1902) );
  NAND2_X1 U489 ( .A1(n1902), .A2(b[4]), .ZN(n118) );
  OAI211_X1 U490 ( .C1(n1448), .C2(n1611), .A(n119), .B(n118), .ZN(n121) );
  NAND2_X1 U491 ( .A1(n1517), .A2(a[19]), .ZN(n1449) );
  NOR2_X1 U492 ( .A1(n1449), .A2(b[5]), .ZN(n120) );
  NOR2_X1 U493 ( .A1(n121), .A2(n120), .ZN(n1239) );
  NAND2_X1 U494 ( .A1(n883), .A2(n125), .ZN(n1722) );
  NOR2_X1 U495 ( .A1(n1722), .A2(b[13]), .ZN(n128) );
  NOR2_X1 U496 ( .A1(n123), .A2(a[11]), .ZN(n1725) );
  NAND2_X1 U497 ( .A1(n1725), .A2(b[12]), .ZN(n122) );
  OAI21_X1 U498 ( .B1(n1702), .B2(b[12]), .A(n122), .ZN(n127) );
  NAND3_X1 U499 ( .A1(n125), .A2(n124), .A3(n123), .ZN(n1723) );
  NOR2_X1 U500 ( .A1(n1723), .A2(n1670), .ZN(n126) );
  NOR3_X1 U501 ( .A1(n128), .A2(n127), .A3(n126), .ZN(n1241) );
  XNOR2_X1 U502 ( .A(n1239), .B(n1241), .ZN(n134) );
  NOR2_X1 U503 ( .A1(n130), .A2(a[19]), .ZN(n1881) );
  INV_X1 U504 ( .A(a[20]), .ZN(n129) );
  NAND2_X1 U505 ( .A1(n1881), .A2(n129), .ZN(n190) );
  NAND2_X1 U506 ( .A1(n158), .A2(n130), .ZN(n1883) );
  MUX2_X1 U507 ( .A(n190), .B(n1883), .S(b[2]), .Z(n133) );
  XNOR2_X1 U508 ( .A(a[19]), .B(a[20]), .ZN(n1391) );
  NOR2_X1 U509 ( .A1(n1391), .A2(a[21]), .ZN(n1374) );
  NAND2_X1 U510 ( .A1(n1374), .A2(b[3]), .ZN(n132) );
  NOR2_X1 U511 ( .A1(n1391), .A2(n130), .ZN(n1884) );
  NAND2_X1 U512 ( .A1(n1884), .A2(n1787), .ZN(n131) );
  NAND3_X1 U513 ( .A1(n133), .A2(n132), .A3(n131), .ZN(n1238) );
  XNOR2_X1 U514 ( .A(n134), .B(n1238), .ZN(n1426) );
  NOR2_X1 U515 ( .A1(a[21]), .A2(a[22]), .ZN(n438) );
  NOR2_X1 U518 ( .A1(n2166), .A2(a[23]), .ZN(n1999) );
  NOR2_X1 U519 ( .A1(n1234), .A2(n438), .ZN(n1231) );
  NAND2_X1 U520 ( .A1(a[23]), .A2(b[0]), .ZN(n1300) );
  XNOR2_X1 U521 ( .A(n1300), .B(b[1]), .ZN(n136) );
  AOI22_X1 U522 ( .A1(n1135), .A2(b[0]), .B1(n1231), .B2(n136), .ZN(n1214) );
  AOI22_X1 U523 ( .A1(b[15]), .A2(n1697), .B1(n1698), .B2(n1131), .ZN(n137) );
  OAI21_X1 U524 ( .B1(n1701), .B2(b[14]), .A(n138), .ZN(n139) );
  AOI21_X1 U525 ( .B1(n1742), .B2(b[14]), .A(n139), .ZN(n1215) );
  XOR2_X1 U526 ( .A(n1214), .B(n1215), .Z(n143) );
  NOR2_X1 U527 ( .A1(n1770), .A2(n893), .ZN(n142) );
  NOR2_X1 U528 ( .A1(n1769), .A2(b[17]), .ZN(n141) );
  MUX2_X1 U529 ( .A(n1712), .B(n1711), .S(b[16]), .Z(n140) );
  NOR3_X1 U530 ( .A1(n142), .A2(n141), .A3(n140), .ZN(n1216) );
  XOR2_X1 U531 ( .A(n143), .B(n1216), .Z(n1423) );
  XNOR2_X1 U532 ( .A(n1426), .B(n1423), .ZN(n174) );
  MUX2_X1 U533 ( .A(n144), .B(n1788), .S(n893), .Z(n146) );
  MUX2_X1 U534 ( .A(n1789), .B(n1599), .S(b[16]), .Z(n145) );
  NAND2_X1 U535 ( .A1(n146), .A2(n145), .ZN(n1446) );
  NOR2_X1 U536 ( .A1(n1770), .A2(n1131), .ZN(n149) );
  NOR2_X1 U537 ( .A1(n1769), .A2(b[15]), .ZN(n148) );
  MUX2_X1 U538 ( .A(n1712), .B(n1711), .S(b[14]), .Z(n147) );
  NOR3_X1 U539 ( .A1(n149), .A2(n148), .A3(n147), .ZN(n1445) );
  NOR2_X1 U542 ( .A1(n627), .A2(n633), .ZN(n1583) );
  NAND3_X1 U543 ( .A1(n633), .A2(a[13]), .A3(a[14]), .ZN(n833) );
  NOR2_X1 U544 ( .A1(a[14]), .A2(n633), .ZN(n831) );
  NAND2_X1 U545 ( .A1(n232), .A2(n831), .ZN(n1481) );
  NOR2_X1 U546 ( .A1(n1481), .A2(b[6]), .ZN(n151) );
  AOI21_X1 U547 ( .B1(n1579), .B2(b[6]), .A(n151), .ZN(n153) );
  NAND2_X1 U548 ( .A1(n1478), .A2(b[7]), .ZN(n152) );
  NAND2_X1 U549 ( .A1(n153), .A2(n152), .ZN(n154) );
  AOI21_X1 U550 ( .B1(n1583), .B2(n1735), .A(n154), .ZN(n1444) );
  NAND2_X1 U551 ( .A1(n1445), .A2(n1444), .ZN(n157) );
  INV_X1 U552 ( .A(n1445), .ZN(n156) );
  INV_X1 U553 ( .A(n1444), .ZN(n155) );
  AOI22_X1 U554 ( .A1(n1446), .A2(n157), .B1(n156), .B2(n155), .ZN(n173) );
  NAND2_X1 U557 ( .A1(n159), .A2(a[21]), .ZN(n2009) );
  NOR2_X1 U560 ( .A1(n173), .A2(n1379), .ZN(n1472) );
  MUX2_X1 U561 ( .A(n1850), .B(n1849), .S(b[19]), .Z(n163) );
  MUX2_X1 U562 ( .A(n1852), .B(n1851), .S(b[18]), .Z(n162) );
  NAND2_X1 U563 ( .A1(n163), .A2(n162), .ZN(n1466) );
  NAND2_X1 U567 ( .A1(n1466), .A2(n1464), .ZN(n172) );
  NOR2_X1 U568 ( .A1(n1722), .A2(b[11]), .ZN(n169) );
  NAND2_X1 U569 ( .A1(n1725), .A2(b[10]), .ZN(n166) );
  OAI21_X1 U570 ( .B1(n1702), .B2(b[10]), .A(n166), .ZN(n168) );
  NOR2_X1 U571 ( .A1(n1723), .A2(n1717), .ZN(n167) );
  NOR3_X1 U572 ( .A1(n169), .A2(n168), .A3(n167), .ZN(n1465) );
  INV_X1 U573 ( .A(n1466), .ZN(n171) );
  INV_X1 U574 ( .A(n1464), .ZN(n170) );
  AOI22_X1 U575 ( .A1(n172), .A2(n1465), .B1(n171), .B2(n170), .ZN(n1475) );
  NAND2_X1 U576 ( .A1(n173), .A2(n1379), .ZN(n1473) );
  OAI21_X1 U577 ( .B1(n1472), .B2(n1475), .A(n1473), .ZN(n1422) );
  XNOR2_X1 U578 ( .A(n174), .B(n1422), .ZN(n368) );
  NAND2_X1 U581 ( .A1(\intadd_79/n1 ), .A2(\intadd_52/SUM[1] ), .ZN(n367) );
  NOR2_X1 U582 ( .A1(n367), .A2(n368), .ZN(n1944) );
  NOR2_X1 U583 ( .A1(\intadd_79/n1 ), .A2(\intadd_52/SUM[1] ), .ZN(n369) );
  NOR2_X1 U584 ( .A1(n177), .A2(n368), .ZN(n178) );
  NOR3_X1 U585 ( .A1(n179), .A2(n1944), .A3(n178), .ZN(n588) );
  XNOR2_X1 U586 ( .A(n180), .B(n588), .ZN(\intadd_57/B[3] ) );
  NOR2_X1 U587 ( .A1(a[12]), .A2(a[11]), .ZN(n649) );
  NAND2_X1 U588 ( .A1(\intadd_69/A[0] ), .A2(n181), .ZN(n1616) );
  NOR2_X1 U589 ( .A1(n1706), .A2(a[13]), .ZN(n1617) );
  AOI21_X1 U592 ( .B1(n1617), .B2(b[23]), .A(n183), .ZN(n184) );
  NAND2_X1 U593 ( .A1(n1616), .A2(n184), .ZN(n239) );
  NAND2_X1 U594 ( .A1(a[23]), .A2(b[12]), .ZN(n238) );
  XNOR2_X1 U595 ( .A(n239), .B(n238), .ZN(n189) );
  NOR2_X1 U596 ( .A1(n1481), .A2(b[21]), .ZN(n185) );
  AOI21_X1 U597 ( .B1(n1579), .B2(b[21]), .A(n185), .ZN(n188) );
  NAND2_X1 U598 ( .A1(n1583), .A2(n1996), .ZN(n187) );
  NAND2_X1 U599 ( .A1(n1478), .A2(b[22]), .ZN(n186) );
  NAND3_X1 U600 ( .A1(n188), .A2(n187), .A3(n186), .ZN(n240) );
  XOR2_X1 U601 ( .A(n189), .B(n240), .Z(n210) );
  NOR2_X1 U602 ( .A1(n1883), .A2(n1602), .ZN(n191) );
  AOI21_X1 U603 ( .B1(n1377), .B2(n1602), .A(n191), .ZN(n194) );
  NAND2_X1 U604 ( .A1(n1884), .A2(n1131), .ZN(n193) );
  NAND2_X1 U605 ( .A1(n1374), .A2(b[15]), .ZN(n192) );
  NAND3_X1 U606 ( .A1(n194), .A2(n193), .A3(n192), .ZN(n881) );
  NOR2_X1 U607 ( .A1(n1481), .A2(b[20]), .ZN(n195) );
  AOI21_X1 U608 ( .B1(n1579), .B2(b[20]), .A(n195), .ZN(n198) );
  NAND2_X1 U609 ( .A1(n1583), .A2(n1991), .ZN(n197) );
  NAND2_X1 U610 ( .A1(n1478), .A2(b[21]), .ZN(n196) );
  NAND3_X1 U611 ( .A1(n198), .A2(n197), .A3(n196), .ZN(n879) );
  AND2_X1 U612 ( .A1(n881), .A2(n879), .ZN(n203) );
  NAND2_X1 U613 ( .A1(n1231), .A2(a[23]), .ZN(n1994) );
  INV_X1 U614 ( .A(n1994), .ZN(n1876) );
  NAND2_X1 U615 ( .A1(n1876), .A2(n1670), .ZN(n202) );
  AND2_X1 U616 ( .A1(n1999), .A2(b[12]), .ZN(n199) );
  AOI21_X1 U617 ( .B1(n1869), .B2(n1273), .A(n199), .ZN(n201) );
  NOR2_X1 U618 ( .A1(n1289), .A2(a[23]), .ZN(n1893) );
  NAND2_X1 U619 ( .A1(n1893), .A2(b[13]), .ZN(n200) );
  NAND3_X1 U620 ( .A1(n202), .A2(n201), .A3(n200), .ZN(n880) );
  OAI22_X1 U621 ( .A1(n203), .A2(n880), .B1(n881), .B2(n879), .ZN(n209) );
  XNOR2_X1 U622 ( .A(n210), .B(n209), .ZN(n204) );
  XNOR2_X1 U623 ( .A(\intadd_81/SUM[0] ), .B(n204), .ZN(\intadd_59/B[3] ) );
  NAND2_X1 U624 ( .A1(\intadd_81/n1 ), .A2(\intadd_69/SUM[2] ), .ZN(n206) );
  NOR2_X1 U625 ( .A1(\intadd_81/n1 ), .A2(\intadd_69/SUM[2] ), .ZN(n205) );
  AOI21_X1 U626 ( .B1(n207), .B2(n206), .A(n205), .ZN(n261) );
  NAND2_X1 U627 ( .A1(\intadd_69/SUM[3] ), .A2(n261), .ZN(n2133) );
  XNOR2_X1 U628 ( .A(\intadd_69/SUM[2] ), .B(\intadd_68/SUM[1] ), .ZN(n208) );
  XNOR2_X1 U629 ( .A(n208), .B(\intadd_81/n1 ), .ZN(n258) );
  NAND2_X1 U630 ( .A1(\intadd_81/SUM[2] ), .A2(\intadd_69/SUM[1] ), .ZN(n256)
         );
  OAI21_X1 U631 ( .B1(\intadd_81/SUM[0] ), .B2(n210), .A(n209), .ZN(n212) );
  NAND2_X1 U632 ( .A1(\intadd_81/SUM[0] ), .A2(n210), .ZN(n211) );
  NAND2_X1 U633 ( .A1(n212), .A2(n211), .ZN(n878) );
  NOR2_X1 U635 ( .A1(a[15]), .A2(a[16]), .ZN(n213) );
  NAND2_X1 U636 ( .A1(n293), .A2(n782), .ZN(n1394) );
  NOR2_X1 U637 ( .A1(n1394), .A2(b[19]), .ZN(n219) );
  NAND2_X1 U639 ( .A1(n1530), .A2(b[18]), .ZN(n217) );
  NOR3_X1 U640 ( .A1(n215), .A2(a[15]), .A3(a[16]), .ZN(n1531) );
  NAND2_X1 U641 ( .A1(n1531), .A2(n1247), .ZN(n216) );
  OAI211_X1 U642 ( .C1(n1437), .C2(n1341), .A(n217), .B(n216), .ZN(n218) );
  NOR2_X1 U646 ( .A1(n1883), .A2(n1131), .ZN(n221) );
  AOI21_X1 U647 ( .B1(n1377), .B2(n1131), .A(n221), .ZN(n224) );
  NAND2_X1 U648 ( .A1(n1884), .A2(n1246), .ZN(n223) );
  NAND2_X1 U649 ( .A1(n1374), .A2(b[16]), .ZN(n222) );
  NAND3_X1 U650 ( .A1(n224), .A2(n223), .A3(n222), .ZN(n251) );
  OAI21_X1 U651 ( .B1(b[10]), .B2(b[11]), .A(a[23]), .ZN(n914) );
  NAND2_X1 U652 ( .A1(n251), .A2(n225), .ZN(n226) );
  NOR2_X1 U653 ( .A1(n253), .A2(n226), .ZN(n909) );
  NAND2_X1 U654 ( .A1(n1902), .A2(b[16]), .ZN(n227) );
  OAI21_X1 U655 ( .B1(n1450), .B2(b[16]), .A(n227), .ZN(n228) );
  AOI21_X1 U656 ( .B1(n989), .B2(b[17]), .A(n228), .ZN(n230) );
  NAND2_X1 U657 ( .A1(n1900), .A2(n893), .ZN(n229) );
  NAND2_X1 U658 ( .A1(n230), .A2(n229), .ZN(n885) );
  INV_X1 U659 ( .A(n885), .ZN(n237) );
  NOR3_X1 U661 ( .A1(n232), .A2(a[11]), .A3(a[12]), .ZN(n1618) );
  AOI22_X1 U662 ( .A1(n1389), .A2(b[23]), .B1(n1618), .B2(n1996), .ZN(n234) );
  NAND2_X1 U663 ( .A1(n1617), .A2(b[22]), .ZN(n233) );
  OAI211_X1 U664 ( .C1(b[23]), .C2(n1616), .A(n234), .B(n233), .ZN(n884) );
  NAND2_X1 U665 ( .A1(n884), .A2(n1730), .ZN(n236) );
  INV_X1 U666 ( .A(n884), .ZN(n235) );
  AOI22_X1 U667 ( .A1(n237), .A2(n236), .B1(n235), .B2(n883), .ZN(n912) );
  AOI21_X1 U668 ( .B1(n240), .B2(n239), .A(n238), .ZN(n242) );
  NOR2_X1 U669 ( .A1(n240), .A2(n239), .ZN(n241) );
  NOR2_X1 U670 ( .A1(n242), .A2(n241), .ZN(n864) );
  NAND2_X1 U671 ( .A1(n1374), .A2(b[17]), .ZN(n244) );
  NAND2_X1 U672 ( .A1(n1377), .A2(n1246), .ZN(n243) );
  OAI211_X1 U673 ( .C1(n1246), .C2(n1883), .A(n244), .B(n243), .ZN(n245) );
  AOI21_X1 U674 ( .B1(n1884), .B2(n893), .A(n245), .ZN(n859) );
  NAND2_X1 U675 ( .A1(n1876), .A2(n1131), .ZN(n249) );
  AND2_X1 U676 ( .A1(n1999), .A2(b[14]), .ZN(n246) );
  AOI21_X1 U677 ( .B1(n1869), .B2(n1602), .A(n246), .ZN(n248) );
  NAND2_X1 U678 ( .A1(n1893), .A2(b[15]), .ZN(n247) );
  NAND3_X1 U679 ( .A1(n249), .A2(n248), .A3(n247), .ZN(n863) );
  XOR2_X1 U680 ( .A(n859), .B(n863), .Z(n250) );
  XNOR2_X1 U681 ( .A(n864), .B(n250), .ZN(n254) );
  OAI21_X1 U682 ( .B1(n253), .B2(n914), .A(n252), .ZN(n910) );
  OAI211_X1 U683 ( .C1(n909), .C2(n912), .A(n254), .B(n910), .ZN(n875) );
  AOI211_X1 U684 ( .C1(n910), .C2(n912), .A(n254), .B(n909), .ZN(n874) );
  AOI21_X1 U685 ( .B1(n878), .B2(n875), .A(n874), .ZN(n259) );
  NOR2_X1 U686 ( .A1(\intadd_81/SUM[2] ), .A2(\intadd_69/SUM[1] ), .ZN(n255)
         );
  AOI21_X1 U687 ( .B1(n256), .B2(n259), .A(n255), .ZN(n257) );
  NAND2_X1 U688 ( .A1(n258), .A2(n257), .ZN(n2130) );
  NAND2_X1 U689 ( .A1(n2133), .A2(n2130), .ZN(n2026) );
  NOR2_X1 U690 ( .A1(n258), .A2(n257), .ZN(n2025) );
  XOR2_X1 U691 ( .A(\intadd_69/SUM[1] ), .B(n259), .Z(n260) );
  XNOR2_X1 U692 ( .A(\intadd_81/SUM[2] ), .B(n260), .ZN(n602) );
  NOR2_X1 U693 ( .A1(\intadd_60/n1 ), .A2(n602), .ZN(n1937) );
  NOR2_X1 U694 ( .A1(n2025), .A2(n1937), .ZN(n2023) );
  NOR2_X1 U695 ( .A1(n2026), .A2(n2023), .ZN(n2033) );
  NOR2_X1 U696 ( .A1(\intadd_69/SUM[3] ), .A2(n261), .ZN(n2032) );
  NOR2_X1 U697 ( .A1(\intadd_69/n1 ), .A2(\intadd_68/SUM[3] ), .ZN(n2027) );
  NOR2_X1 U698 ( .A1(n2032), .A2(n2027), .ZN(n2138) );
  INV_X1 U699 ( .A(n2138), .ZN(n262) );
  NOR2_X1 U700 ( .A1(n2033), .A2(n262), .ZN(n2146) );
  NAND2_X1 U701 ( .A1(\intadd_69/n1 ), .A2(\intadd_68/SUM[3] ), .ZN(n2036) );
  NAND2_X1 U702 ( .A1(n1439), .A2(n1996), .ZN(n264) );
  NAND2_X1 U703 ( .A1(n1902), .A2(b[22]), .ZN(n263) );
  OAI211_X1 U704 ( .C1(n1448), .C2(n2165), .A(n264), .B(n263), .ZN(n266) );
  NOR2_X1 U705 ( .A1(n1449), .A2(b[23]), .ZN(n265) );
  NOR2_X1 U706 ( .A1(n266), .A2(n265), .ZN(n301) );
  OAI21_X1 U708 ( .B1(b[17]), .B2(b[16]), .A(a[23]), .ZN(n267) );
  AOI21_X1 U709 ( .B1(n301), .B2(n268), .A(n267), .ZN(n309) );
  NAND2_X1 U710 ( .A1(n1876), .A2(n1309), .ZN(n272) );
  AND2_X1 U711 ( .A1(n1999), .A2(b[19]), .ZN(n269) );
  AOI21_X1 U712 ( .B1(n1869), .B2(n1341), .A(n269), .ZN(n271) );
  NAND2_X1 U713 ( .A1(n1893), .A2(b[20]), .ZN(n270) );
  NAND3_X1 U714 ( .A1(n272), .A2(n271), .A3(n270), .ZN(n307) );
  XNOR2_X1 U715 ( .A(n309), .B(n307), .ZN(n284) );
  NAND2_X1 U716 ( .A1(n1893), .A2(b[19]), .ZN(n275) );
  NAND2_X1 U717 ( .A1(n1999), .A2(b[18]), .ZN(n274) );
  NAND2_X1 U718 ( .A1(n1869), .A2(n1247), .ZN(n273) );
  NAND3_X1 U719 ( .A1(n275), .A2(n274), .A3(n273), .ZN(n277) );
  NOR2_X1 U720 ( .A1(n1994), .A2(b[19]), .ZN(n276) );
  NOR2_X1 U721 ( .A1(n277), .A2(n276), .ZN(n285) );
  NOR2_X1 U722 ( .A1(n1883), .A2(n1309), .ZN(n278) );
  AOI21_X1 U723 ( .B1(n1377), .B2(n1309), .A(n278), .ZN(n281) );
  NAND2_X1 U724 ( .A1(n1884), .A2(n1991), .ZN(n280) );
  NAND2_X1 U725 ( .A1(n1374), .A2(b[21]), .ZN(n279) );
  NAND3_X1 U726 ( .A1(n281), .A2(n280), .A3(n279), .ZN(n287) );
  NAND2_X1 U727 ( .A1(n287), .A2(n770), .ZN(n283) );
  NOR2_X1 U728 ( .A1(n287), .A2(n770), .ZN(n282) );
  AOI21_X1 U729 ( .B1(n285), .B2(n283), .A(n282), .ZN(n308) );
  XNOR2_X1 U730 ( .A(n284), .B(n308), .ZN(n321) );
  XNOR2_X1 U731 ( .A(\intadd_58/SUM[0] ), .B(n321), .ZN(n305) );
  INV_X1 U732 ( .A(n285), .ZN(n286) );
  XNOR2_X1 U733 ( .A(n286), .B(n770), .ZN(n288) );
  XNOR2_X1 U734 ( .A(n288), .B(n287), .ZN(n820) );
  NAND2_X1 U735 ( .A1(n1902), .A2(b[21]), .ZN(n289) );
  OAI21_X1 U736 ( .B1(n1450), .B2(b[21]), .A(n289), .ZN(n290) );
  AOI21_X1 U737 ( .B1(n989), .B2(b[22]), .A(n290), .ZN(n292) );
  NAND2_X1 U738 ( .A1(n1900), .A2(n1996), .ZN(n291) );
  NAND2_X1 U739 ( .A1(n292), .A2(n291), .ZN(n809) );
  NAND2_X1 U740 ( .A1(n1530), .A2(b[23]), .ZN(n295) );
  NAND2_X1 U741 ( .A1(n293), .A2(n2165), .ZN(n294) );
  NAND3_X1 U742 ( .A1(n1394), .A2(n295), .A3(n294), .ZN(n808) );
  NAND2_X1 U743 ( .A1(n809), .A2(n808), .ZN(n298) );
  AND2_X1 U744 ( .A1(a[23]), .A2(b[16]), .ZN(n807) );
  INV_X1 U745 ( .A(n809), .ZN(n297) );
  AOI22_X1 U746 ( .A1(n298), .A2(n807), .B1(n297), .B2(n296), .ZN(n817) );
  NAND2_X1 U747 ( .A1(n820), .A2(n817), .ZN(n304) );
  XNOR2_X1 U750 ( .A(n301), .B(n300), .ZN(n818) );
  INV_X1 U751 ( .A(n820), .ZN(n303) );
  INV_X1 U752 ( .A(n817), .ZN(n302) );
  AOI22_X1 U753 ( .A1(n304), .A2(n818), .B1(n303), .B2(n302), .ZN(n324) );
  XNOR2_X1 U754 ( .A(n305), .B(n324), .ZN(n306) );
  NAND2_X1 U755 ( .A1(\intadd_68/n1 ), .A2(n306), .ZN(n2039) );
  NAND2_X1 U756 ( .A1(n2036), .A2(n2039), .ZN(n2137) );
  NOR2_X1 U757 ( .A1(\intadd_68/n1 ), .A2(n306), .ZN(n2140) );
  NAND2_X1 U759 ( .A1(n308), .A2(n309), .ZN(n312) );
  NOR2_X1 U762 ( .A1(n1883), .A2(n1996), .ZN(n314) );
  AOI21_X1 U763 ( .B1(n1377), .B2(n1996), .A(n314), .ZN(n317) );
  NAND2_X1 U764 ( .A1(n1884), .A2(n2165), .ZN(n316) );
  NAND2_X1 U765 ( .A1(n1374), .A2(b[23]), .ZN(n315) );
  NAND3_X1 U766 ( .A1(n317), .A2(n316), .A3(n315), .ZN(n654) );
  XNOR2_X1 U769 ( .A(n654), .B(n319), .ZN(n607) );
  XOR2_X1 U770 ( .A(n326), .B(n607), .Z(n320) );
  XNOR2_X1 U771 ( .A(\intadd_58/SUM[1] ), .B(n320), .ZN(n331) );
  INV_X1 U772 ( .A(n331), .ZN(n325) );
  INV_X1 U773 ( .A(n321), .ZN(n322) );
  NAND2_X1 U774 ( .A1(\intadd_58/SUM[0] ), .A2(n322), .ZN(n323) );
  OAI21_X1 U775 ( .B1(n2), .B2(n324), .A(n323), .ZN(n329) );
  NOR2_X1 U776 ( .A1(n325), .A2(n329), .ZN(n2142) );
  AOI21_X1 U777 ( .B1(n2037), .B2(n2150), .A(n2149), .ZN(n610) );
  NAND2_X1 U778 ( .A1(\intadd_58/SUM[1] ), .A2(n327), .ZN(n605) );
  NOR2_X1 U779 ( .A1(\intadd_58/SUM[1] ), .A2(n327), .ZN(n608) );
  AOI21_X1 U780 ( .B1(n605), .B2(n607), .A(n608), .ZN(n328) );
  NAND2_X1 U781 ( .A1(\intadd_58/SUM[2] ), .A2(n328), .ZN(n2153) );
  INV_X1 U782 ( .A(n329), .ZN(n330) );
  NOR2_X1 U783 ( .A1(n331), .A2(n330), .ZN(n2152) );
  INV_X1 U784 ( .A(n2152), .ZN(n332) );
  NAND2_X1 U785 ( .A1(n2153), .A2(n332), .ZN(n2154) );
  AOI22_X1 U786 ( .A1(\intadd_46/n2 ), .A2(n334), .B1(n333), .B2(
        \intadd_46/A[4] ), .ZN(n335) );
  NAND2_X1 U787 ( .A1(\intadd_66/SUM[2] ), .A2(\intadd_75/n1 ), .ZN(n339) );
  NOR2_X1 U788 ( .A1(n339), .A2(n341), .ZN(n340) );
  NOR2_X1 U790 ( .A1(\intadd_66/SUM[2] ), .A2(\intadd_75/n1 ), .ZN(n346) );
  AOI21_X1 U791 ( .B1(n339), .B2(n341), .A(n346), .ZN(n345) );
  NAND2_X1 U792 ( .A1(\intadd_66/SUM[3] ), .A2(n345), .ZN(n2094) );
  AOI21_X1 U793 ( .B1(n346), .B2(\intadd_65/SUM[1] ), .A(n340), .ZN(n344) );
  NAND2_X1 U796 ( .A1(n344), .A2(n343), .ZN(n2060) );
  NAND2_X1 U797 ( .A1(n2060), .A2(\intadd_64/n1 ), .ZN(n2057) );
  NAND2_X1 U798 ( .A1(n2094), .A2(n2057), .ZN(n350) );
  NOR2_X1 U799 ( .A1(\intadd_66/SUM[3] ), .A2(n345), .ZN(n2093) );
  NOR3_X1 U800 ( .A1(\intadd_64/n1 ), .A2(\intadd_65/SUM[1] ), .A3(n347), .ZN(
        n348) );
  NOR2_X1 U801 ( .A1(n2093), .A2(n348), .ZN(n349) );
  OAI21_X1 U802 ( .B1(n351), .B2(n350), .A(n349), .ZN(n1907) );
  NAND2_X1 U803 ( .A1(\intadd_65/SUM[3] ), .A2(\intadd_66/n1 ), .ZN(n1905) );
  NAND2_X1 U804 ( .A1(\intadd_76/SUM[2] ), .A2(n1903), .ZN(n1979) );
  NAND2_X1 U805 ( .A1(n1979), .A2(n1904), .ZN(n352) );
  AOI21_X1 U806 ( .B1(n1907), .B2(n1905), .A(n352), .ZN(n1912) );
  NAND2_X1 U807 ( .A1(n1912), .A2(n1982), .ZN(n366) );
  NAND2_X1 U808 ( .A1(\intadd_55/SUM[4] ), .A2(\intadd_57/A[1] ), .ZN(n354) );
  NAND2_X1 U809 ( .A1(\intadd_77/SUM[2] ), .A2(n353), .ZN(n1981) );
  OAI211_X1 U810 ( .C1(n1913), .C2(n1910), .A(n354), .B(n1981), .ZN(n355) );
  AOI21_X1 U811 ( .B1(\intadd_77/n1 ), .B2(\intadd_57/B[0] ), .A(n355), .ZN(
        n365) );
  NAND2_X1 U812 ( .A1(n357), .A2(n356), .ZN(n358) );
  OAI22_X1 U813 ( .A1(\intadd_56/SUM[4] ), .A2(\intadd_55/n1 ), .B1(
        \intadd_77/n1 ), .B2(n358), .ZN(n363) );
  NAND2_X1 U814 ( .A1(n360), .A2(n359), .ZN(n361) );
  AOI21_X1 U815 ( .B1(n361), .B2(\intadd_57/A[1] ), .A(\intadd_55/SUM[4] ), 
        .ZN(n362) );
  AOI21_X1 U816 ( .B1(n366), .B2(n365), .A(n364), .ZN(n379) );
  OAI21_X1 U817 ( .B1(n369), .B2(n368), .A(n367), .ZN(n569) );
  XOR2_X1 U818 ( .A(n569), .B(\intadd_52/SUM[2] ), .Z(n370) );
  XNOR2_X1 U819 ( .A(\intadd_53/SUM[3] ), .B(n370), .ZN(n2063) );
  OAI21_X1 U820 ( .B1(n1942), .B2(n588), .A(n371), .ZN(n2062) );
  AOI22_X1 U821 ( .A1(\intadd_57/B[3] ), .A2(\intadd_56/n1 ), .B1(
        \intadd_55/n1 ), .B2(\intadd_56/SUM[4] ), .ZN(n372) );
  OAI21_X1 U822 ( .B1(n2063), .B2(n373), .A(n372), .ZN(n378) );
  AOI22_X1 U823 ( .A1(\intadd_56/n1 ), .A2(n2062), .B1(n375), .B2(n374), .ZN(
        n376) );
  NAND2_X1 U824 ( .A1(n2063), .A2(n376), .ZN(n377) );
  OAI21_X1 U825 ( .B1(n379), .B2(n378), .A(n377), .ZN(n1947) );
  NAND2_X1 U826 ( .A1(\intadd_50/SUM[3] ), .A2(\intadd_71/SUM[2] ), .ZN(n580)
         );
  NOR2_X1 U829 ( .A1(n382), .A2(n581), .ZN(n383) );
  XNOR2_X1 U830 ( .A(n383), .B(n582), .ZN(n591) );
  NAND2_X1 U831 ( .A1(\intadd_63/SUM[3] ), .A2(\intadd_61/n1 ), .ZN(n410) );
  NOR2_X1 U832 ( .A1(n1722), .A2(b[19]), .ZN(n387) );
  NAND2_X1 U833 ( .A1(n1725), .A2(b[18]), .ZN(n384) );
  OAI21_X1 U834 ( .B1(n1702), .B2(b[18]), .A(n384), .ZN(n386) );
  NOR2_X1 U835 ( .A1(n1723), .A2(n1341), .ZN(n385) );
  NOR3_X1 U836 ( .A1(n387), .A2(n386), .A3(n385), .ZN(n1080) );
  NOR2_X1 U837 ( .A1(n1394), .A2(b[13]), .ZN(n391) );
  NAND2_X1 U838 ( .A1(n1530), .A2(b[12]), .ZN(n389) );
  NAND2_X1 U839 ( .A1(n1531), .A2(n1273), .ZN(n388) );
  OAI211_X1 U840 ( .C1(n1437), .C2(n1670), .A(n389), .B(n388), .ZN(n390) );
  NOR2_X1 U841 ( .A1(n391), .A2(n390), .ZN(n1079) );
  XNOR2_X1 U842 ( .A(n1080), .B(n1079), .ZN(n395) );
  MUX2_X1 U843 ( .A(n1698), .B(n1697), .S(b[21]), .Z(n394) );
  NOR2_X1 U844 ( .A1(n1701), .A2(b[20]), .ZN(n392) );
  AOI21_X1 U845 ( .B1(b[20]), .B2(n1742), .A(n392), .ZN(n393) );
  NAND2_X1 U846 ( .A1(n394), .A2(n393), .ZN(n1083) );
  XNOR2_X1 U847 ( .A(n395), .B(n1083), .ZN(n1123) );
  AOI22_X1 U848 ( .A1(b[16]), .A2(n1617), .B1(n1618), .B2(n1246), .ZN(n396) );
  OAI21_X1 U849 ( .B1(n1619), .B2(n893), .A(n396), .ZN(n397) );
  INV_X1 U850 ( .A(n397), .ZN(n398) );
  OAI21_X1 U851 ( .B1(b[17]), .B2(n1616), .A(n398), .ZN(n400) );
  NAND2_X1 U852 ( .A1(a[23]), .A2(b[4]), .ZN(n1136) );
  NAND2_X1 U853 ( .A1(a[23]), .A2(b[5]), .ZN(n399) );
  NAND2_X1 U854 ( .A1(n1136), .A2(n399), .ZN(n401) );
  INV_X1 U855 ( .A(n1136), .ZN(n1092) );
  NAND2_X1 U856 ( .A1(n1092), .A2(b[5]), .ZN(n1066) );
  NAND2_X1 U857 ( .A1(n1066), .A2(n401), .ZN(n402) );
  AOI22_X1 U858 ( .A1(n1068), .A2(n1066), .B1(n403), .B2(n402), .ZN(n1122) );
  INV_X1 U859 ( .A(n1122), .ZN(n405) );
  AOI22_X1 U860 ( .A1(n406), .A2(n405), .B1(n404), .B2(\intadd_71/SUM[0] ), 
        .ZN(n1098) );
  XOR2_X1 U861 ( .A(\intadd_49/SUM[1] ), .B(n1098), .Z(n407) );
  XNOR2_X1 U862 ( .A(n407), .B(\intadd_71/SUM[1] ), .ZN(n411) );
  INV_X1 U863 ( .A(n411), .ZN(n409) );
  NOR2_X1 U864 ( .A1(\intadd_63/SUM[3] ), .A2(\intadd_61/n1 ), .ZN(n408) );
  AOI21_X1 U865 ( .B1(n410), .B2(n409), .A(n408), .ZN(n590) );
  NAND2_X1 U866 ( .A1(n591), .A2(n590), .ZN(n2103) );
  XNOR2_X1 U867 ( .A(\intadd_61/n1 ), .B(n411), .ZN(n412) );
  XNOR2_X1 U868 ( .A(n412), .B(\intadd_63/SUM[3] ), .ZN(n1954) );
  NAND2_X1 U869 ( .A1(\intadd_51/n1 ), .A2(n1954), .ZN(n2018) );
  NAND2_X1 U870 ( .A1(n2103), .A2(n2018), .ZN(n2105) );
  NAND2_X1 U872 ( .A1(\intadd_52/SUM[4] ), .A2(\intadd_53/n1 ), .ZN(n2068) );
  NOR2_X1 U873 ( .A1(n1394), .A2(b[10]), .ZN(n417) );
  NAND2_X1 U874 ( .A1(n1530), .A2(b[9]), .ZN(n415) );
  NAND2_X1 U875 ( .A1(n1531), .A2(n1684), .ZN(n414) );
  OAI211_X1 U876 ( .C1(n1732), .C2(n1437), .A(n415), .B(n414), .ZN(n416) );
  NOR2_X1 U877 ( .A1(n417), .A2(n416), .ZN(n449) );
  AOI22_X1 U878 ( .A1(b[16]), .A2(n1723), .B1(n1722), .B2(n1246), .ZN(n418) );
  AOI21_X1 U879 ( .B1(n1725), .B2(b[15]), .A(n418), .ZN(n419) );
  OAI21_X1 U880 ( .B1(n1702), .B2(b[15]), .A(n419), .ZN(n450) );
  XNOR2_X1 U881 ( .A(n449), .B(n450), .ZN(n423) );
  AOI22_X1 U882 ( .A1(b[11]), .A2(n833), .B1(n1481), .B2(n1717), .ZN(n420) );
  AOI21_X1 U883 ( .B1(n1478), .B2(b[12]), .A(n420), .ZN(n422) );
  NAND2_X1 U884 ( .A1(n1583), .A2(n1273), .ZN(n421) );
  NAND2_X1 U885 ( .A1(n422), .A2(n421), .ZN(n452) );
  XNOR2_X1 U886 ( .A(n423), .B(n452), .ZN(n523) );
  NAND2_X1 U887 ( .A1(n1439), .A2(n1735), .ZN(n425) );
  NAND2_X1 U888 ( .A1(n1902), .A2(b[7]), .ZN(n424) );
  OAI211_X1 U889 ( .C1(n1448), .C2(n1694), .A(n425), .B(n424), .ZN(n427) );
  NOR2_X1 U890 ( .A1(n1449), .A2(b[8]), .ZN(n426) );
  NOR2_X1 U891 ( .A1(n427), .A2(n426), .ZN(n458) );
  INV_X1 U892 ( .A(n1557), .ZN(n1506) );
  NAND3_X1 U893 ( .A1(a[7]), .A2(b[17]), .A3(n1250), .ZN(n428) );
  NAND2_X1 U894 ( .A1(n1506), .A2(n428), .ZN(n431) );
  XNOR2_X1 U895 ( .A(a[9]), .B(b[18]), .ZN(n429) );
  NAND2_X1 U896 ( .A1(n1666), .A2(n429), .ZN(n430) );
  AOI22_X1 U897 ( .A1(n431), .A2(n430), .B1(n1741), .B2(n893), .ZN(n456) );
  XNOR2_X1 U898 ( .A(n458), .B(n456), .ZN(n435) );
  NOR2_X1 U899 ( .A1(n1770), .A2(n1309), .ZN(n434) );
  NOR2_X1 U900 ( .A1(n1769), .A2(b[20]), .ZN(n433) );
  MUX2_X1 U901 ( .A(n1712), .B(n1711), .S(b[19]), .Z(n432) );
  NOR3_X1 U902 ( .A1(n434), .A2(n433), .A3(n432), .ZN(n457) );
  OAI21_X1 U904 ( .B1(\intadd_61/SUM[0] ), .B2(n523), .A(n525), .ZN(n437) );
  NAND2_X1 U905 ( .A1(\intadd_61/SUM[0] ), .A2(n523), .ZN(n436) );
  NAND2_X1 U906 ( .A1(n437), .A2(n436), .ZN(n1194) );
  NOR2_X1 U907 ( .A1(n1994), .A2(b[3]), .ZN(n1189) );
  NAND2_X1 U908 ( .A1(n1189), .A2(n1611), .ZN(n443) );
  AOI22_X1 U909 ( .A1(n1893), .A2(b[5]), .B1(b[4]), .B2(n1999), .ZN(n442) );
  AND2_X1 U910 ( .A1(n1869), .A2(n1651), .ZN(n440) );
  AND2_X1 U911 ( .A1(a[23]), .A2(b[3]), .ZN(n1138) );
  AOI22_X1 U912 ( .A1(n1231), .A2(n1611), .B1(n438), .B2(n1651), .ZN(n439) );
  OAI22_X1 U913 ( .A1(n440), .A2(n1138), .B1(n439), .B2(n1787), .ZN(n441) );
  NAND3_X1 U914 ( .A1(n443), .A2(n442), .A3(n441), .ZN(n447) );
  AOI22_X1 U915 ( .A1(b[15]), .A2(n1619), .B1(n1616), .B2(n1131), .ZN(n444) );
  AOI21_X1 U916 ( .B1(n1618), .B2(n1602), .A(n444), .ZN(n446) );
  NAND2_X1 U917 ( .A1(n1617), .A2(b[14]), .ZN(n445) );
  NAND2_X1 U918 ( .A1(n446), .A2(n445), .ZN(n1137) );
  XNOR2_X1 U919 ( .A(n447), .B(n1137), .ZN(n1165) );
  NOR2_X1 U920 ( .A1(n449), .A2(n448), .ZN(n453) );
  INV_X1 U921 ( .A(n449), .ZN(n451) );
  OAI22_X1 U922 ( .A1(n453), .A2(n452), .B1(n451), .B2(n450), .ZN(n1167) );
  XNOR2_X1 U923 ( .A(n1165), .B(n1167), .ZN(n460) );
  AOI22_X1 U926 ( .A1(n459), .A2(n458), .B1(n457), .B2(n456), .ZN(n1170) );
  XOR2_X1 U927 ( .A(n460), .B(n1170), .Z(n1193) );
  XNOR2_X1 U928 ( .A(n1194), .B(n1193), .ZN(n477) );
  NOR2_X1 U929 ( .A1(n1770), .A2(n1991), .ZN(n463) );
  NOR2_X1 U930 ( .A1(n1769), .A2(b[21]), .ZN(n462) );
  MUX2_X1 U931 ( .A(n1712), .B(n1711), .S(b[20]), .Z(n461) );
  NOR3_X1 U932 ( .A1(n463), .A2(n462), .A3(n461), .ZN(n1114) );
  NOR2_X1 U933 ( .A1(n1883), .A2(n1859), .ZN(n464) );
  AOI21_X1 U934 ( .B1(n1377), .B2(n1859), .A(n464), .ZN(n467) );
  NAND2_X1 U935 ( .A1(n1884), .A2(n1735), .ZN(n466) );
  NAND2_X1 U936 ( .A1(n1374), .A2(b[7]), .ZN(n465) );
  NAND3_X1 U937 ( .A1(n467), .A2(n466), .A3(n465), .ZN(n1119) );
  XNOR2_X1 U938 ( .A(n1114), .B(n1119), .ZN(n470) );
  MUX2_X1 U939 ( .A(n144), .B(n1788), .S(n2165), .Z(n469) );
  MUX2_X1 U940 ( .A(n1789), .B(n1599), .S(b[22]), .Z(n468) );
  NAND2_X1 U941 ( .A1(n469), .A2(n468), .ZN(n1118) );
  XNOR2_X1 U942 ( .A(n470), .B(n1118), .ZN(n534) );
  NOR2_X1 U943 ( .A1(n1481), .A2(b[12]), .ZN(n471) );
  AOI21_X1 U944 ( .B1(n1579), .B2(b[12]), .A(n471), .ZN(n474) );
  NAND2_X1 U945 ( .A1(n1583), .A2(n1670), .ZN(n473) );
  NAND2_X1 U946 ( .A1(n1478), .A2(b[13]), .ZN(n472) );
  NAND3_X1 U947 ( .A1(n474), .A2(n473), .A3(n472), .ZN(n1147) );
  NAND3_X1 U948 ( .A1(n475), .A2(a[3]), .A3(a[1]), .ZN(n1172) );
  NAND2_X1 U949 ( .A1(n1331), .A2(n1205), .ZN(n1174) );
  NAND2_X1 U950 ( .A1(n1172), .A2(n1174), .ZN(n509) );
  XNOR2_X1 U951 ( .A(n1147), .B(n509), .ZN(n532) );
  XNOR2_X1 U952 ( .A(n534), .B(n532), .ZN(n476) );
  XNOR2_X1 U953 ( .A(\intadd_63/SUM[0] ), .B(n476), .ZN(n1197) );
  XOR2_X1 U954 ( .A(n477), .B(n1197), .Z(n563) );
  XNOR2_X1 U955 ( .A(\intadd_62/n1 ), .B(n563), .ZN(n528) );
  NAND2_X1 U956 ( .A1(n1439), .A2(n1859), .ZN(n479) );
  NAND2_X1 U957 ( .A1(n1902), .A2(b[6]), .ZN(n478) );
  OAI211_X1 U958 ( .C1(n1448), .C2(n1735), .A(n479), .B(n478), .ZN(n481) );
  NOR2_X1 U959 ( .A1(n1449), .A2(b[7]), .ZN(n480) );
  NOR2_X1 U960 ( .A1(n481), .A2(n480), .ZN(n520) );
  AOI22_X1 U961 ( .A1(b[17]), .A2(n1697), .B1(n1698), .B2(n893), .ZN(n482) );
  OAI21_X1 U962 ( .B1(n1701), .B2(b[16]), .A(n483), .ZN(n484) );
  AOI21_X1 U963 ( .B1(n1742), .B2(b[16]), .A(n484), .ZN(n518) );
  XNOR2_X1 U964 ( .A(n520), .B(n518), .ZN(n488) );
  NOR2_X1 U965 ( .A1(n1770), .A2(n1341), .ZN(n487) );
  NOR2_X1 U966 ( .A1(n1769), .A2(b[19]), .ZN(n486) );
  MUX2_X1 U967 ( .A(n1712), .B(n1711), .S(b[18]), .Z(n485) );
  NOR3_X1 U968 ( .A1(n487), .A2(n486), .A3(n485), .ZN(n519) );
  XNOR2_X1 U969 ( .A(n488), .B(n519), .ZN(n1345) );
  NOR2_X1 U970 ( .A1(n1394), .A2(b[9]), .ZN(n492) );
  NAND2_X1 U971 ( .A1(n1530), .A2(b[8]), .ZN(n490) );
  NAND2_X1 U972 ( .A1(n1531), .A2(n1694), .ZN(n489) );
  OAI211_X1 U973 ( .C1(n1684), .C2(n1437), .A(n490), .B(n489), .ZN(n491) );
  NOR2_X1 U974 ( .A1(n492), .A2(n491), .ZN(n502) );
  AOI22_X1 U975 ( .A1(b[15]), .A2(n1723), .B1(n1722), .B2(n1131), .ZN(n493) );
  AOI21_X1 U976 ( .B1(n1725), .B2(b[14]), .A(n493), .ZN(n494) );
  OAI21_X1 U977 ( .B1(n1702), .B2(b[14]), .A(n494), .ZN(n504) );
  XOR2_X1 U978 ( .A(n502), .B(n504), .Z(n499) );
  NOR2_X1 U979 ( .A1(n1481), .A2(b[10]), .ZN(n495) );
  AOI21_X1 U980 ( .B1(n1579), .B2(b[10]), .A(n495), .ZN(n497) );
  NAND2_X1 U981 ( .A1(n1478), .A2(b[11]), .ZN(n496) );
  NAND2_X1 U982 ( .A1(n497), .A2(n496), .ZN(n498) );
  AOI21_X1 U983 ( .B1(n1583), .B2(n1717), .A(n498), .ZN(n503) );
  XNOR2_X1 U984 ( .A(n499), .B(n503), .ZN(n1344) );
  OAI21_X1 U985 ( .B1(\intadd_51/SUM[0] ), .B2(n1345), .A(n1344), .ZN(n501) );
  NAND2_X1 U986 ( .A1(\intadd_51/SUM[0] ), .A2(n1345), .ZN(n500) );
  NAND2_X1 U987 ( .A1(n501), .A2(n500), .ZN(n1212) );
  INV_X1 U988 ( .A(n502), .ZN(n506) );
  INV_X1 U989 ( .A(n503), .ZN(n505) );
  AOI21_X1 U990 ( .B1(n506), .B2(n505), .A(n504), .ZN(n508) );
  NOR2_X1 U991 ( .A1(n506), .A2(n505), .ZN(n507) );
  NOR2_X1 U992 ( .A1(n508), .A2(n507), .ZN(n1199) );
  NOR2_X1 U993 ( .A1(n1171), .A2(n1327), .ZN(n513) );
  NAND2_X1 U994 ( .A1(a[23]), .A2(b[2]), .ZN(n1186) );
  AOI21_X1 U995 ( .B1(n513), .B2(n1172), .A(n1186), .ZN(n511) );
  INV_X1 U996 ( .A(n509), .ZN(n512) );
  NAND2_X1 U997 ( .A1(n512), .A2(n2165), .ZN(n510) );
  NAND2_X1 U998 ( .A1(n511), .A2(n510), .ZN(n515) );
  OAI211_X1 U999 ( .C1(n513), .C2(n2165), .A(n512), .B(n1186), .ZN(n514) );
  NAND2_X1 U1000 ( .A1(n515), .A2(n514), .ZN(n1201) );
  XNOR2_X1 U1001 ( .A(n1199), .B(n1201), .ZN(n522) );
  AOI22_X1 U1005 ( .A1(n521), .A2(n520), .B1(n519), .B2(n518), .ZN(n1200) );
  XOR2_X1 U1006 ( .A(n522), .B(n1200), .Z(n1210) );
  XOR2_X1 U1008 ( .A(\intadd_61/SUM[0] ), .B(n526), .Z(n1211) );
  FA_X1 U1009 ( .A(n1212), .B(n1210), .CI(n1211), .CO(n529), .S() );
  XNOR2_X1 U1010 ( .A(\intadd_73/n1 ), .B(n529), .ZN(n527) );
  XNOR2_X1 U1011 ( .A(n527), .B(\intadd_51/SUM[2] ), .ZN(n564) );
  XNOR2_X1 U1012 ( .A(n528), .B(n564), .ZN(n574) );
  NAND2_X1 U1013 ( .A1(\intadd_52/n1 ), .A2(n574), .ZN(n2070) );
  OAI21_X1 U1014 ( .B1(\intadd_51/SUM[2] ), .B2(\intadd_73/n1 ), .A(n529), 
        .ZN(n531) );
  NAND2_X1 U1015 ( .A1(\intadd_51/SUM[2] ), .A2(\intadd_73/n1 ), .ZN(n530) );
  NAND2_X1 U1016 ( .A1(n531), .A2(n530), .ZN(n558) );
  INV_X1 U1017 ( .A(n532), .ZN(n533) );
  OAI21_X1 U1018 ( .B1(\intadd_63/SUM[0] ), .B2(n534), .A(n533), .ZN(n536) );
  NAND2_X1 U1019 ( .A1(\intadd_63/SUM[0] ), .A2(n534), .ZN(n535) );
  NAND2_X1 U1020 ( .A1(n536), .A2(n535), .ZN(n1160) );
  XNOR2_X1 U1021 ( .A(\intadd_63/SUM[1] ), .B(n1160), .ZN(n556) );
  NAND2_X1 U1022 ( .A1(n1876), .A2(n1859), .ZN(n540) );
  AND2_X1 U1023 ( .A1(n1999), .A2(b[5]), .ZN(n537) );
  AOI21_X1 U1024 ( .B1(n1869), .B2(n1611), .A(n537), .ZN(n539) );
  NAND2_X1 U1025 ( .A1(n1893), .A2(b[6]), .ZN(n538) );
  NAND3_X1 U1026 ( .A1(n540), .A2(n539), .A3(n538), .ZN(n1108) );
  NOR2_X1 U1027 ( .A1(n1722), .A2(b[18]), .ZN(n544) );
  NAND2_X1 U1028 ( .A1(n1725), .A2(b[17]), .ZN(n541) );
  OAI21_X1 U1029 ( .B1(n1702), .B2(b[17]), .A(n541), .ZN(n543) );
  NOR2_X1 U1030 ( .A1(n1723), .A2(n1247), .ZN(n542) );
  NOR3_X1 U1031 ( .A1(n544), .A2(n543), .A3(n542), .ZN(n1107) );
  XNOR2_X1 U1032 ( .A(n1108), .B(n1107), .ZN(n548) );
  MUX2_X1 U1033 ( .A(n1698), .B(n1697), .S(b[20]), .Z(n547) );
  NOR2_X1 U1034 ( .A1(n1701), .A2(b[19]), .ZN(n545) );
  AOI21_X1 U1035 ( .B1(b[19]), .B2(n1742), .A(n545), .ZN(n546) );
  NAND2_X1 U1036 ( .A1(n547), .A2(n546), .ZN(n1110) );
  XNOR2_X1 U1037 ( .A(n548), .B(n1110), .ZN(n1125) );
  NAND2_X1 U1038 ( .A1(n1331), .A2(a[5]), .ZN(n549) );
  MUX2_X1 U1039 ( .A(n549), .B(n1599), .S(b[23]), .Z(n550) );
  NAND2_X1 U1040 ( .A1(n550), .A2(n1788), .ZN(n1095) );
  XOR2_X1 U1041 ( .A(n1095), .B(n1136), .Z(n554) );
  NOR2_X1 U1042 ( .A1(n1770), .A2(n1996), .ZN(n553) );
  NOR2_X1 U1043 ( .A1(n1769), .A2(b[22]), .ZN(n552) );
  MUX2_X1 U1044 ( .A(n1712), .B(n1711), .S(b[21]), .Z(n551) );
  NOR3_X1 U1045 ( .A1(n553), .A2(n552), .A3(n551), .ZN(n1091) );
  XOR2_X1 U1046 ( .A(n554), .B(n1091), .Z(n1126) );
  XNOR2_X1 U1047 ( .A(n1125), .B(n1126), .ZN(n555) );
  XOR2_X1 U1048 ( .A(\intadd_50/SUM[0] ), .B(n555), .Z(n1161) );
  XOR2_X1 U1049 ( .A(n556), .B(n1161), .Z(n557) );
  NAND2_X1 U1050 ( .A1(\intadd_51/SUM[3] ), .A2(n561), .ZN(n559) );
  NAND2_X1 U1051 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U1052 ( .A1(n559), .A2(n560), .ZN(n577) );
  NAND2_X1 U1053 ( .A1(\intadd_51/SUM[4] ), .A2(n577), .ZN(n1966) );
  NAND2_X1 U1054 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U1055 ( .A(\intadd_51/SUM[3] ), .B(n562), .Z(n573) );
  NAND3_X1 U1059 ( .A1(n586), .A2(n1952), .A3(n2016), .ZN(n1919) );
  NAND2_X1 U1062 ( .A1(\intadd_53/SUM[4] ), .A2(n1949), .ZN(n1917) );
  NOR2_X1 U1064 ( .A1(\intadd_53/SUM[4] ), .A2(n1949), .ZN(n576) );
  NAND2_X1 U1065 ( .A1(n573), .A2(n572), .ZN(n1953) );
  INV_X1 U1066 ( .A(n1953), .ZN(n2098) );
  NOR2_X1 U1067 ( .A1(\intadd_52/SUM[4] ), .A2(\intadd_53/n1 ), .ZN(n2069) );
  NAND2_X1 U1068 ( .A1(n2069), .A2(n2070), .ZN(n575) );
  NAND2_X1 U1069 ( .A1(n575), .A2(n2071), .ZN(n1951) );
  AOI211_X1 U1070 ( .C1(n1952), .C2(n576), .A(n2098), .B(n1951), .ZN(n579) );
  NOR2_X1 U1071 ( .A1(\intadd_51/SUM[4] ), .A2(n577), .ZN(n1965) );
  NOR2_X1 U1072 ( .A1(\intadd_51/n1 ), .A2(n1954), .ZN(n2019) );
  NOR2_X1 U1073 ( .A1(n1965), .A2(n2019), .ZN(n2107) );
  OAI21_X1 U1074 ( .B1(n579), .B2(n578), .A(n2107), .ZN(n587) );
  OAI21_X1 U1075 ( .B1(n582), .B2(n581), .A(n580), .ZN(n583) );
  NOR2_X1 U1076 ( .A1(\intadd_50/SUM[4] ), .A2(n583), .ZN(n1960) );
  NOR2_X1 U1077 ( .A1(\intadd_50/n1 ), .A2(\intadd_49/SUM[4] ), .ZN(n2079) );
  NOR2_X1 U1078 ( .A1(n1960), .A2(n2079), .ZN(n2112) );
  NOR2_X1 U1079 ( .A1(\intadd_49/n1 ), .A2(\intadd_47/SUM[4] ), .ZN(n2114) );
  INV_X1 U1080 ( .A(n2114), .ZN(n584) );
  OAI21_X1 U1081 ( .B1(n2112), .B2(n2111), .A(n584), .ZN(n585) );
  AOI21_X1 U1082 ( .B1(n587), .B2(n586), .A(n585), .ZN(n1925) );
  NAND2_X1 U1083 ( .A1(n1942), .A2(n588), .ZN(n589) );
  NOR2_X1 U1084 ( .A1(\intadd_56/n1 ), .A2(n589), .ZN(n1915) );
  NOR2_X1 U1085 ( .A1(n591), .A2(n590), .ZN(n2106) );
  NOR2_X1 U1086 ( .A1(n2111), .A2(n2104), .ZN(n1921) );
  AOI22_X1 U1087 ( .A1(n593), .A2(n592), .B1(n1921), .B2(n2076), .ZN(n594) );
  NOR2_X1 U1089 ( .A1(\intadd_48/SUM[4] ), .A2(\intadd_47/n1 ), .ZN(n1987) );
  NOR2_X1 U1090 ( .A1(\intadd_48/n1 ), .A2(\intadd_59/SUM[3] ), .ZN(n2122) );
  NOR2_X1 U1091 ( .A1(\intadd_59/n1 ), .A2(\intadd_60/SUM[3] ), .ZN(n597) );
  NOR3_X1 U1092 ( .A1(n1987), .A2(n2122), .A3(n597), .ZN(n1924) );
  NOR2_X1 U1093 ( .A1(n2115), .A2(n1988), .ZN(n1933) );
  NAND2_X1 U1094 ( .A1(\intadd_59/A[3] ), .A2(\intadd_59/B[3] ), .ZN(n598) );
  NAND2_X1 U1095 ( .A1(n2118), .A2(n598), .ZN(n599) );
  AOI22_X1 U1096 ( .A1(n2125), .A2(n599), .B1(\intadd_60/SUM[3] ), .B2(
        \intadd_59/n1 ), .ZN(n1916) );
  AOI21_X1 U1097 ( .B1(n601), .B2(n1924), .A(n600), .ZN(n1927) );
  NAND2_X1 U1098 ( .A1(n602), .A2(\intadd_60/n1 ), .ZN(n2024) );
  INV_X1 U1099 ( .A(n2024), .ZN(n1930) );
  NOR3_X1 U1100 ( .A1(n2029), .A2(n2137), .A3(n2154), .ZN(n603) );
  OAI211_X1 U1101 ( .C1(n1986), .C2(n604), .A(n1927), .B(n603), .ZN(n609) );
  INV_X1 U1102 ( .A(\intadd_58/SUM[2] ), .ZN(n606) );
  OAI211_X1 U1103 ( .C1(n608), .C2(n607), .A(n606), .B(n605), .ZN(n2157) );
  OAI211_X1 U1104 ( .C1(n610), .C2(n2154), .A(n609), .B(n2157), .ZN(n611) );
  AOI22_X1 U1105 ( .A1(b[17]), .A2(n1478), .B1(n1583), .B2(n893), .ZN(n612) );
  OAI21_X1 U1106 ( .B1(n1481), .B2(b[16]), .A(n612), .ZN(n613) );
  AOI21_X1 U1107 ( .B1(n1579), .B2(b[16]), .A(n613), .ZN(n618) );
  NOR2_X1 U1110 ( .A1(n618), .A2(n615), .ZN(n1002) );
  NAND2_X1 U1111 ( .A1(b[6]), .A2(b[7]), .ZN(n619) );
  NAND2_X1 U1112 ( .A1(n616), .A2(n619), .ZN(n617) );
  AOI22_X1 U1113 ( .A1(n1002), .A2(n619), .B1(n618), .B2(n617), .ZN(n620) );
  INV_X2 U1114 ( .A(\intadd_53/SUM[1] ), .ZN(\intadd_78/B[2] ) );
  INV_X2 U1115 ( .A(\intadd_77/SUM[1] ), .ZN(\intadd_76/B[2] ) );
  INV_X2 U1116 ( .A(\intadd_67/SUM[2] ), .ZN(\intadd_76/A[2] ) );
  INV_X2 U1117 ( .A(\intadd_76/SUM[1] ), .ZN(\intadd_65/B[3] ) );
  INV_X2 U1118 ( .A(\intadd_67/SUM[1] ), .ZN(\intadd_76/A[1] ) );
  MUX2_X1 U1119 ( .A(n1619), .B(n1616), .S(n1740), .Z(n622) );
  MUX2_X1 U1120 ( .A(n1596), .B(n1276), .S(b[1]), .Z(n621) );
  NOR2_X1 U1121 ( .A1(n1722), .A2(b[4]), .ZN(n626) );
  NAND2_X1 U1122 ( .A1(n1725), .A2(b[3]), .ZN(n623) );
  OAI21_X1 U1123 ( .B1(n1702), .B2(b[3]), .A(n623), .ZN(n625) );
  NOR2_X1 U1124 ( .A1(n1723), .A2(n1651), .ZN(n624) );
  NOR3_X1 U1125 ( .A1(n626), .A2(n625), .A3(n624), .ZN(n1646) );
  NAND2_X1 U1126 ( .A1(n628), .A2(n1646), .ZN(n630) );
  NOR2_X1 U1127 ( .A1(n627), .A2(n2084), .ZN(n1645) );
  INV_X1 U1128 ( .A(n1646), .ZN(n629) );
  AOI22_X1 U1129 ( .A1(n630), .A2(n1645), .B1(n629), .B2(n1647), .ZN(n1674) );
  MUX2_X1 U1130 ( .A(n1850), .B(n1849), .S(b[13]), .Z(n632) );
  MUX2_X1 U1131 ( .A(n1852), .B(n1851), .S(b[12]), .Z(n631) );
  NAND2_X1 U1132 ( .A1(n632), .A2(n631), .ZN(n1672) );
  AND2_X1 U1133 ( .A1(n1478), .A2(b[1]), .ZN(n637) );
  AOI21_X1 U1134 ( .B1(a[13]), .B2(a[14]), .A(n633), .ZN(n844) );
  OAI21_X1 U1135 ( .B1(n2086), .B2(n2084), .A(n844), .ZN(n634) );
  OAI211_X1 U1136 ( .C1(n833), .C2(n2084), .A(n1481), .B(n634), .ZN(n636) );
  NAND2_X1 U1137 ( .A1(n2084), .A2(n844), .ZN(n635) );
  AOI21_X1 U1138 ( .B1(n1481), .B2(b[1]), .A(n635), .ZN(n1627) );
  OAI21_X1 U1139 ( .B1(n637), .B2(n636), .A(n1629), .ZN(n1671) );
  INV_X1 U1140 ( .A(n1671), .ZN(n638) );
  NAND2_X1 U1141 ( .A1(n1672), .A2(n638), .ZN(n640) );
  AOI22_X1 U1142 ( .A1(n1674), .A2(n640), .B1(n639), .B2(n1671), .ZN(n641) );
  INV_X2 U1143 ( .A(\intadd_67/SUM[0] ), .ZN(\intadd_76/CI ) );
  INV_X2 U1144 ( .A(\intadd_54/n1 ), .ZN(\intadd_46/B[3] ) );
  OAI21_X1 U1145 ( .B1(n643), .B2(n642), .A(n1799), .ZN(n644) );
  INV_X1 U1146 ( .A(n644), .ZN(\intadd_72/B[0] ) );
  NAND2_X1 U1147 ( .A1(n1062), .A2(n2086), .ZN(n646) );
  AOI21_X1 U1148 ( .B1(n646), .B2(n1752), .A(b[0]), .ZN(\intadd_54/A[0] ) );
  INV_X2 U1149 ( .A(\intadd_46/SUM[2] ), .ZN(\intadd_54/A[4] ) );
  INV_X2 U1150 ( .A(\intadd_74/SUM[2] ), .ZN(\intadd_46/A[3] ) );
  INV_X2 U1151 ( .A(\intadd_64/SUM[2] ), .ZN(\intadd_74/B[2] ) );
  INV_X2 U1152 ( .A(\intadd_75/SUM[1] ), .ZN(\intadd_74/A[2] ) );
  MUX2_X1 U1153 ( .A(n1619), .B(n1616), .S(n2086), .Z(n648) );
  MUX2_X1 U1154 ( .A(n1596), .B(n1276), .S(b[0]), .Z(n647) );
  NOR2_X1 U1155 ( .A1(n2084), .A2(n649), .ZN(n1707) );
  NAND2_X1 U1156 ( .A1(\intadd_69/A[0] ), .A2(n650), .ZN(n651) );
  NOR2_X1 U1157 ( .A1(n652), .A2(n651), .ZN(n1692) );
  AOI21_X1 U1158 ( .B1(n652), .B2(n651), .A(n1692), .ZN(n653) );
  INV_X2 U1159 ( .A(n653), .ZN(\intadd_75/A[1] ) );
  AOI21_X1 U1160 ( .B1(b[19]), .B2(b[18]), .A(n654), .ZN(n655) );
  AOI211_X1 U1161 ( .C1(n1341), .C2(n1247), .A(n2167), .B(n655), .ZN(n656) );
  INV_X1 U1162 ( .A(n656), .ZN(\intadd_58/B[2] ) );
  MUX2_X1 U1163 ( .A(n1531), .B(n1530), .S(b[20]), .Z(n657) );
  AOI21_X1 U1164 ( .B1(b[21]), .B2(n1529), .A(n657), .ZN(n658) );
  OAI21_X1 U1165 ( .B1(b[21]), .B2(n1394), .A(n658), .ZN(n867) );
  AOI21_X1 U1166 ( .B1(b[12]), .B2(b[13]), .A(n867), .ZN(n659) );
  AOI211_X1 U1167 ( .C1(n1670), .C2(n1273), .A(n2167), .B(n659), .ZN(n660) );
  INV_X1 U1168 ( .A(n660), .ZN(\intadd_69/B[1] ) );
  NOR2_X1 U1169 ( .A1(n1883), .A2(n1670), .ZN(n661) );
  AOI21_X1 U1170 ( .B1(n1377), .B2(n1670), .A(n661), .ZN(n664) );
  NAND2_X1 U1171 ( .A1(n1884), .A2(n1602), .ZN(n663) );
  NAND2_X1 U1172 ( .A1(n1374), .A2(b[14]), .ZN(n662) );
  AND3_X1 U1173 ( .A1(n664), .A2(n663), .A3(n662), .ZN(n2182) );
  NOR2_X1 U1174 ( .A1(n1883), .A2(n1694), .ZN(n665) );
  AOI21_X1 U1175 ( .B1(n1377), .B2(n1694), .A(n665), .ZN(n668) );
  NAND2_X1 U1176 ( .A1(n1884), .A2(n1684), .ZN(n667) );
  NAND2_X1 U1177 ( .A1(n1374), .A2(b[9]), .ZN(n666) );
  AND3_X1 U1178 ( .A1(n668), .A2(n667), .A3(n666), .ZN(n2183) );
  NOR2_X1 U1179 ( .A1(n1883), .A2(n1651), .ZN(n669) );
  AOI21_X1 U1180 ( .B1(n1377), .B2(n1651), .A(n669), .ZN(n672) );
  NAND2_X1 U1181 ( .A1(n1884), .A2(n1611), .ZN(n671) );
  NAND2_X1 U1182 ( .A1(n1374), .A2(b[5]), .ZN(n670) );
  AND3_X1 U1183 ( .A1(n672), .A2(n671), .A3(n670), .ZN(n2184) );
  NOR2_X1 U1184 ( .A1(n1883), .A2(n1735), .ZN(n673) );
  AOI21_X1 U1185 ( .B1(n1377), .B2(n1735), .A(n673), .ZN(n676) );
  NAND2_X1 U1186 ( .A1(n1884), .A2(n1694), .ZN(n675) );
  NAND2_X1 U1187 ( .A1(n1374), .A2(b[8]), .ZN(n674) );
  AND3_X1 U1188 ( .A1(n676), .A2(n675), .A3(n674), .ZN(n2185) );
  NOR2_X1 U1189 ( .A1(n1883), .A2(n1611), .ZN(n677) );
  AOI21_X1 U1190 ( .B1(n1377), .B2(n1611), .A(n677), .ZN(n680) );
  NAND2_X1 U1191 ( .A1(n1884), .A2(n1859), .ZN(n679) );
  NAND2_X1 U1192 ( .A1(n1374), .A2(b[6]), .ZN(n678) );
  AND3_X1 U1193 ( .A1(n680), .A2(n679), .A3(n678), .ZN(n2186) );
  NOR2_X1 U1194 ( .A1(n1883), .A2(n893), .ZN(n681) );
  AOI21_X1 U1195 ( .B1(n1377), .B2(n893), .A(n681), .ZN(n684) );
  NAND2_X1 U1196 ( .A1(n1884), .A2(n1247), .ZN(n683) );
  NAND2_X1 U1197 ( .A1(n1374), .A2(b[18]), .ZN(n682) );
  AND3_X1 U1198 ( .A1(n684), .A2(n683), .A3(n682), .ZN(n2187) );
  NOR2_X1 U1199 ( .A1(n1481), .A2(b[22]), .ZN(n685) );
  AOI21_X1 U1200 ( .B1(n1579), .B2(b[22]), .A(n685), .ZN(n688) );
  NAND2_X1 U1201 ( .A1(n1583), .A2(n2165), .ZN(n687) );
  NAND2_X1 U1202 ( .A1(n1478), .A2(b[23]), .ZN(n686) );
  AND3_X1 U1203 ( .A1(n688), .A2(n687), .A3(n686), .ZN(n2188) );
  NOR2_X1 U1204 ( .A1(n1481), .A2(b[3]), .ZN(n689) );
  AOI21_X1 U1205 ( .B1(n1579), .B2(b[3]), .A(n689), .ZN(n692) );
  NAND2_X1 U1206 ( .A1(n1583), .A2(n1651), .ZN(n691) );
  NAND2_X1 U1207 ( .A1(n1478), .A2(b[4]), .ZN(n690) );
  AND3_X1 U1208 ( .A1(n692), .A2(n691), .A3(n690), .ZN(n2189) );
  NOR2_X1 U1209 ( .A1(n1481), .A2(b[15]), .ZN(n693) );
  AOI21_X1 U1210 ( .B1(n1579), .B2(b[15]), .A(n693), .ZN(n696) );
  NAND2_X1 U1211 ( .A1(n1583), .A2(n1246), .ZN(n695) );
  NAND2_X1 U1212 ( .A1(n1478), .A2(b[16]), .ZN(n694) );
  AND3_X1 U1213 ( .A1(n696), .A2(n695), .A3(n694), .ZN(n2190) );
  NOR2_X1 U1214 ( .A1(n1883), .A2(n1991), .ZN(n697) );
  AOI21_X1 U1215 ( .B1(n1377), .B2(n1991), .A(n697), .ZN(n700) );
  NAND2_X1 U1216 ( .A1(n1884), .A2(n1996), .ZN(n699) );
  NAND2_X1 U1217 ( .A1(n1374), .A2(b[22]), .ZN(n698) );
  AND3_X1 U1218 ( .A1(n700), .A2(n699), .A3(n698), .ZN(n2191) );
  NOR2_X1 U1219 ( .A1(n1883), .A2(n1684), .ZN(n701) );
  AOI21_X1 U1220 ( .B1(n1377), .B2(n1684), .A(n701), .ZN(n704) );
  NAND2_X1 U1221 ( .A1(n1884), .A2(n1732), .ZN(n703) );
  NAND2_X1 U1222 ( .A1(n1374), .A2(b[10]), .ZN(n702) );
  AND3_X1 U1223 ( .A1(n704), .A2(n703), .A3(n702), .ZN(n2192) );
  NOR2_X1 U1224 ( .A1(n1481), .A2(b[14]), .ZN(n705) );
  AOI21_X1 U1225 ( .B1(n1579), .B2(b[14]), .A(n705), .ZN(n708) );
  NAND2_X1 U1226 ( .A1(n1583), .A2(n1131), .ZN(n707) );
  NAND2_X1 U1227 ( .A1(n1478), .A2(b[15]), .ZN(n706) );
  AND3_X1 U1228 ( .A1(n708), .A2(n707), .A3(n706), .ZN(n2193) );
  NOR2_X1 U1229 ( .A1(n1883), .A2(n1732), .ZN(n709) );
  AOI21_X1 U1230 ( .B1(n1377), .B2(n1732), .A(n709), .ZN(n712) );
  NAND2_X1 U1231 ( .A1(n1884), .A2(n1717), .ZN(n711) );
  NAND2_X1 U1232 ( .A1(n1374), .A2(b[11]), .ZN(n710) );
  AND3_X1 U1233 ( .A1(n712), .A2(n711), .A3(n710), .ZN(n2194) );
  NOR2_X1 U1234 ( .A1(n1883), .A2(n1273), .ZN(n713) );
  AOI21_X1 U1235 ( .B1(n1377), .B2(n1273), .A(n713), .ZN(n716) );
  NAND2_X1 U1236 ( .A1(n1884), .A2(n1670), .ZN(n715) );
  NAND2_X1 U1237 ( .A1(n1374), .A2(b[13]), .ZN(n714) );
  AND3_X1 U1238 ( .A1(n716), .A2(n715), .A3(n714), .ZN(n2195) );
  NOR2_X1 U1239 ( .A1(n1481), .A2(b[8]), .ZN(n717) );
  AOI21_X1 U1240 ( .B1(n1579), .B2(b[8]), .A(n717), .ZN(n720) );
  NAND2_X1 U1241 ( .A1(n1583), .A2(n1684), .ZN(n719) );
  NAND2_X1 U1242 ( .A1(n1478), .A2(b[9]), .ZN(n718) );
  AND3_X1 U1243 ( .A1(n720), .A2(n719), .A3(n718), .ZN(n2196) );
  NOR2_X1 U1244 ( .A1(n1481), .A2(b[19]), .ZN(n721) );
  AOI21_X1 U1245 ( .B1(n1579), .B2(b[19]), .A(n721), .ZN(n724) );
  NAND2_X1 U1246 ( .A1(n1583), .A2(n1309), .ZN(n723) );
  NAND2_X1 U1247 ( .A1(n1478), .A2(b[20]), .ZN(n722) );
  AND3_X1 U1248 ( .A1(n724), .A2(n723), .A3(n722), .ZN(n2197) );
  NOR2_X1 U1249 ( .A1(n1481), .A2(b[7]), .ZN(n725) );
  AOI21_X1 U1250 ( .B1(n1579), .B2(b[7]), .A(n725), .ZN(n728) );
  NAND2_X1 U1251 ( .A1(n1583), .A2(n1694), .ZN(n727) );
  NAND2_X1 U1252 ( .A1(n1478), .A2(b[8]), .ZN(n726) );
  AND3_X1 U1253 ( .A1(n728), .A2(n727), .A3(n726), .ZN(n2198) );
  AOI22_X1 U1254 ( .A1(n1389), .A2(b[7]), .B1(n1618), .B2(n1859), .ZN(n730) );
  NAND2_X1 U1255 ( .A1(n1617), .A2(b[6]), .ZN(n729) );
  OAI211_X1 U1256 ( .C1(b[7]), .C2(n1616), .A(n730), .B(n729), .ZN(n736) );
  NOR2_X1 U1262 ( .A1(n736), .A2(n735), .ZN(n1414) );
  NOR2_X1 U1263 ( .A1(n1395), .A2(n1414), .ZN(n739) );
  NOR2_X1 U1264 ( .A1(n1711), .A2(n1712), .ZN(n1772) );
  XNOR2_X1 U1265 ( .A(a[7]), .B(b[12]), .ZN(n1509) );
  OAI22_X1 U1266 ( .A1(n1770), .A2(n1670), .B1(n1772), .B2(n1509), .ZN(n738)
         );
  NOR2_X1 U1267 ( .A1(n1769), .A2(b[13]), .ZN(n737) );
  NOR2_X1 U1268 ( .A1(n738), .A2(n737), .ZN(n1415) );
  XOR2_X1 U1269 ( .A(n739), .B(n1415), .Z(n1518) );
  AOI22_X1 U1270 ( .A1(n1389), .A2(b[6]), .B1(n1618), .B2(n1611), .ZN(n741) );
  NAND2_X1 U1271 ( .A1(n1617), .A2(b[5]), .ZN(n740) );
  OAI211_X1 U1272 ( .C1(b[6]), .C2(n1616), .A(n741), .B(n740), .ZN(n1535) );
  NAND2_X1 U1276 ( .A1(n1535), .A2(n1534), .ZN(n750) );
  NOR2_X1 U1277 ( .A1(n1722), .A2(b[8]), .ZN(n747) );
  NAND2_X1 U1278 ( .A1(n1725), .A2(b[7]), .ZN(n744) );
  OAI21_X1 U1279 ( .B1(n1702), .B2(b[7]), .A(n744), .ZN(n746) );
  NOR2_X1 U1280 ( .A1(n1723), .A2(n1694), .ZN(n745) );
  NOR3_X1 U1281 ( .A1(n747), .A2(n746), .A3(n745), .ZN(n1536) );
  INV_X1 U1282 ( .A(n1534), .ZN(n749) );
  INV_X1 U1283 ( .A(n1535), .ZN(n748) );
  AOI22_X1 U1284 ( .A1(n750), .A2(n1536), .B1(n749), .B2(n748), .ZN(n1523) );
  XNOR2_X1 U1285 ( .A(n1518), .B(n1523), .ZN(n767) );
  MUX2_X1 U1286 ( .A(n144), .B(n1788), .S(n1131), .Z(n752) );
  MUX2_X1 U1287 ( .A(n1789), .B(n1599), .S(b[14]), .Z(n751) );
  MUX2_X1 U1288 ( .A(n1850), .B(n1849), .S(b[17]), .Z(n754) );
  MUX2_X1 U1289 ( .A(n1852), .B(n1851), .S(b[16]), .Z(n753) );
  NOR2_X1 U1290 ( .A1(n1722), .A2(b[9]), .ZN(n758) );
  NAND2_X1 U1291 ( .A1(n1725), .A2(b[8]), .ZN(n755) );
  OAI21_X1 U1292 ( .B1(n1702), .B2(b[8]), .A(n755), .ZN(n757) );
  NOR2_X1 U1293 ( .A1(n1723), .A2(n1684), .ZN(n756) );
  NOR3_X1 U1294 ( .A1(n758), .A2(n757), .A3(n756), .ZN(n760) );
  NAND2_X1 U1295 ( .A1(n759), .A2(n760), .ZN(n763) );
  INV_X1 U1296 ( .A(n760), .ZN(n761) );
  NAND2_X1 U1297 ( .A1(n762), .A2(n761), .ZN(n1396) );
  NAND2_X1 U1298 ( .A1(n763), .A2(n1396), .ZN(n765) );
  INV_X1 U1299 ( .A(n763), .ZN(n764) );
  NOR2_X1 U1300 ( .A1(n764), .A2(n766), .ZN(n1398) );
  AOI22_X1 U1301 ( .A1(n766), .A2(n765), .B1(n1398), .B2(n1396), .ZN(n1522) );
  XNOR2_X1 U1302 ( .A(n767), .B(n1522), .ZN(\intadd_67/A[3] ) );
  MUX2_X1 U1303 ( .A(n1437), .B(n1394), .S(n2086), .Z(n769) );
  MUX2_X1 U1304 ( .A(n1435), .B(n1434), .S(b[0]), .Z(n768) );
  NAND2_X1 U1305 ( .A1(n769), .A2(n768), .ZN(n772) );
  AOI21_X1 U1306 ( .B1(b[0]), .B2(n1435), .A(n770), .ZN(n771) );
  NAND2_X1 U1307 ( .A1(n772), .A2(n771), .ZN(n1585) );
  NOR2_X1 U1308 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U1309 ( .A1(n1587), .A2(n773), .ZN(n1635) );
  MUX2_X1 U1310 ( .A(n144), .B(n1788), .S(n1670), .Z(n775) );
  MUX2_X1 U1311 ( .A(n1789), .B(n1599), .S(b[12]), .Z(n774) );
  NAND2_X1 U1312 ( .A1(n775), .A2(n774), .ZN(n1633) );
  XNOR2_X1 U1314 ( .A(a[7]), .B(b[11]), .ZN(n1511) );
  NOR2_X1 U1317 ( .A1(n779), .A2(n1632), .ZN(n781) );
  OAI22_X1 U1318 ( .A1(n1635), .A2(n781), .B1(n780), .B2(n1633), .ZN(
        \intadd_67/A[2] ) );
  NAND3_X1 U1319 ( .A1(n783), .A2(b[0]), .A3(n782), .ZN(n1636) );
  INV_X1 U1320 ( .A(n1636), .ZN(n790) );
  OAI22_X1 U1321 ( .A1(n1596), .A2(b[3]), .B1(n1619), .B2(n1651), .ZN(n784) );
  AOI21_X1 U1322 ( .B1(n1617), .B2(b[3]), .A(n784), .ZN(n785) );
  OAI21_X1 U1323 ( .B1(b[4]), .B2(n1616), .A(n785), .ZN(n1637) );
  MUX2_X1 U1324 ( .A(n1583), .B(n1478), .S(b[2]), .Z(n787) );
  MUX2_X1 U1325 ( .A(n1580), .B(n1579), .S(b[1]), .Z(n786) );
  NOR2_X1 U1326 ( .A1(n787), .A2(n786), .ZN(n1638) );
  OAI21_X1 U1327 ( .B1(n788), .B2(n1636), .A(n1638), .ZN(n789) );
  OAI21_X1 U1328 ( .B1(n790), .B2(n1637), .A(n789), .ZN(\intadd_67/A[1] ) );
  MUX2_X1 U1329 ( .A(n1764), .B(n1763), .S(b[14]), .Z(n792) );
  MUX2_X1 U1330 ( .A(n1766), .B(n1765), .S(b[13]), .Z(n791) );
  NOR2_X1 U1331 ( .A1(n792), .A2(n791), .ZN(\intadd_67/A[0] ) );
  NAND2_X1 U1332 ( .A1(n1439), .A2(n1309), .ZN(n794) );
  NAND2_X1 U1333 ( .A1(n1902), .A2(b[20]), .ZN(n793) );
  OAI211_X1 U1334 ( .C1(n1448), .C2(n1991), .A(n794), .B(n793), .ZN(n796) );
  NOR2_X1 U1335 ( .A1(n1449), .A2(b[21]), .ZN(n795) );
  NOR2_X1 U1336 ( .A1(n796), .A2(n795), .ZN(n854) );
  NAND2_X1 U1337 ( .A1(b[15]), .A2(b[14]), .ZN(n797) );
  OAI21_X1 U1338 ( .B1(b[15]), .B2(b[14]), .A(a[23]), .ZN(n852) );
  AOI21_X1 U1339 ( .B1(n854), .B2(n797), .A(n852), .ZN(n842) );
  NOR2_X1 U1340 ( .A1(n1883), .A2(n1341), .ZN(n798) );
  AOI21_X1 U1341 ( .B1(n1377), .B2(n1341), .A(n798), .ZN(n801) );
  NAND2_X1 U1342 ( .A1(n1884), .A2(n1309), .ZN(n800) );
  NAND2_X1 U1343 ( .A1(n1374), .A2(b[20]), .ZN(n799) );
  NAND3_X1 U1344 ( .A1(n801), .A2(n800), .A3(n799), .ZN(n840) );
  INV_X1 U1345 ( .A(n842), .ZN(n805) );
  INV_X1 U1346 ( .A(n840), .ZN(n804) );
  NOR2_X1 U1347 ( .A1(n1994), .A2(b[18]), .ZN(n803) );
  MUX2_X1 U1348 ( .A(n1999), .B(n1869), .S(n893), .Z(n802) );
  AOI211_X1 U1349 ( .C1(n1893), .C2(b[18]), .A(n803), .B(n802), .ZN(n841) );
  OAI21_X1 U1350 ( .B1(n805), .B2(n804), .A(n841), .ZN(n806) );
  OAI21_X1 U1351 ( .B1(n842), .B2(n840), .A(n806), .ZN(\intadd_68/A[3] ) );
  XOR2_X1 U1352 ( .A(n808), .B(n807), .Z(n810) );
  XOR2_X1 U1353 ( .A(n810), .B(n809), .Z(\intadd_68/A[2] ) );
  MUX2_X1 U1354 ( .A(n1435), .B(n1434), .S(b[22]), .Z(n811) );
  OAI21_X1 U1355 ( .B1(n1437), .B2(n2165), .A(n811), .ZN(n812) );
  AOI21_X1 U1356 ( .B1(n1528), .B2(n2165), .A(n812), .ZN(\intadd_68/A[1] ) );
  AND2_X1 U1357 ( .A1(n1893), .A2(b[16]), .ZN(n816) );
  NOR2_X1 U1358 ( .A1(n1994), .A2(b[16]), .ZN(n815) );
  NAND2_X1 U1359 ( .A1(n1999), .A2(b[15]), .ZN(n813) );
  OAI21_X1 U1360 ( .B1(n1895), .B2(b[15]), .A(n813), .ZN(n814) );
  NOR3_X1 U1361 ( .A1(n816), .A2(n815), .A3(n814), .ZN(\intadd_68/A[0] ) );
  XNOR2_X1 U1362 ( .A(n818), .B(n817), .ZN(n819) );
  XNOR2_X1 U1363 ( .A(n820), .B(n819), .ZN(\intadd_68/B[3] ) );
  NAND2_X1 U1364 ( .A1(n1374), .A2(b[19]), .ZN(n822) );
  NAND2_X1 U1365 ( .A1(n1377), .A2(n1247), .ZN(n821) );
  OAI211_X1 U1366 ( .C1(n1883), .C2(n1247), .A(n822), .B(n821), .ZN(n823) );
  AOI21_X1 U1367 ( .B1(n1884), .B2(n1341), .A(n823), .ZN(n846) );
  INV_X1 U1368 ( .A(n846), .ZN(n828) );
  NOR2_X1 U1369 ( .A1(n1994), .A2(b[17]), .ZN(n825) );
  MUX2_X1 U1370 ( .A(n1999), .B(n1869), .S(n1246), .Z(n824) );
  AOI211_X1 U1371 ( .C1(n1893), .C2(b[17]), .A(n825), .B(n824), .ZN(n845) );
  OAI21_X1 U1372 ( .B1(n846), .B2(n844), .A(n845), .ZN(n826) );
  OAI21_X1 U1373 ( .B1(n828), .B2(n827), .A(n826), .ZN(\intadd_68/B[2] ) );
  NAND2_X1 U1374 ( .A1(a[23]), .A2(b[14]), .ZN(n848) );
  MUX2_X1 U1375 ( .A(n1531), .B(n1530), .S(b[21]), .Z(n829) );
  AOI21_X1 U1376 ( .B1(n1529), .B2(b[22]), .A(n829), .ZN(n830) );
  OAI21_X1 U1377 ( .B1(b[22]), .B2(n1394), .A(n830), .ZN(n851) );
  INV_X1 U1378 ( .A(n851), .ZN(n836) );
  NAND2_X1 U1379 ( .A1(n2165), .A2(n831), .ZN(n832) );
  OAI21_X1 U1380 ( .B1(n833), .B2(n2165), .A(n832), .ZN(n834) );
  NOR2_X1 U1381 ( .A1(n1583), .A2(n834), .ZN(n849) );
  OAI21_X1 U1382 ( .B1(n836), .B2(n835), .A(n849), .ZN(n837) );
  OAI21_X1 U1383 ( .B1(n848), .B2(n851), .A(n837), .ZN(\intadd_68/B[1] ) );
  MUX2_X1 U1384 ( .A(n1262), .B(n1450), .S(n1341), .Z(n838) );
  OAI21_X1 U1385 ( .B1(n1309), .B2(n1448), .A(n838), .ZN(n839) );
  AOI21_X1 U1386 ( .B1(n1900), .B2(n1309), .A(n839), .ZN(\intadd_68/CI ) );
  XNOR2_X1 U1387 ( .A(n841), .B(n840), .ZN(n843) );
  XNOR2_X1 U1388 ( .A(n843), .B(n842), .ZN(\intadd_69/A[3] ) );
  XNOR2_X1 U1389 ( .A(n845), .B(n844), .ZN(n847) );
  XNOR2_X1 U1390 ( .A(n847), .B(n846), .ZN(\intadd_69/A[2] ) );
  XOR2_X1 U1391 ( .A(n849), .B(n848), .Z(n850) );
  XOR2_X1 U1392 ( .A(n851), .B(n850), .Z(\intadd_69/A[1] ) );
  AOI21_X1 U1393 ( .B1(b[14]), .B2(b[15]), .A(n852), .ZN(n853) );
  XOR2_X1 U1394 ( .A(n854), .B(n853), .Z(\intadd_69/B[2] ) );
  MUX2_X1 U1395 ( .A(n1262), .B(n1450), .S(n1247), .Z(n855) );
  OAI21_X1 U1396 ( .B1(n1341), .B2(n1448), .A(n855), .ZN(n856) );
  AOI21_X1 U1397 ( .B1(n1900), .B2(n1341), .A(n856), .ZN(\intadd_69/CI ) );
  MUX2_X1 U1398 ( .A(n1435), .B(n1434), .S(b[19]), .Z(n857) );
  OAI21_X1 U1399 ( .B1(n1309), .B2(n1437), .A(n857), .ZN(n858) );
  AOI21_X1 U1400 ( .B1(n1528), .B2(n1309), .A(n858), .ZN(\intadd_81/A[0] ) );
  INV_X1 U1401 ( .A(n864), .ZN(n861) );
  INV_X1 U1402 ( .A(n863), .ZN(n860) );
  OAI21_X1 U1403 ( .B1(n861), .B2(n860), .A(n859), .ZN(n862) );
  OAI21_X1 U1404 ( .B1(n864), .B2(n863), .A(n862), .ZN(\intadd_81/B[2] ) );
  XOR2_X1 U1407 ( .A(n867), .B(n866), .Z(\intadd_81/B[1] ) );
  MUX2_X1 U1408 ( .A(n1262), .B(n1450), .S(n893), .Z(n868) );
  OAI21_X1 U1409 ( .B1(n1247), .B2(n1448), .A(n868), .ZN(n869) );
  AOI21_X1 U1410 ( .B1(n1900), .B2(n1247), .A(n869), .ZN(\intadd_81/B[0] ) );
  AND2_X1 U1411 ( .A1(n1893), .A2(b[14]), .ZN(n873) );
  NOR2_X1 U1412 ( .A1(n1994), .A2(b[14]), .ZN(n872) );
  NAND2_X1 U1413 ( .A1(n1999), .A2(b[13]), .ZN(n870) );
  OAI21_X1 U1414 ( .B1(n1895), .B2(b[13]), .A(n870), .ZN(n871) );
  NOR3_X1 U1415 ( .A1(n873), .A2(n872), .A3(n871), .ZN(\intadd_81/CI ) );
  INV_X1 U1416 ( .A(n874), .ZN(n876) );
  NAND2_X1 U1417 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U1418 ( .A(n878), .B(n877), .ZN(\intadd_60/A[3] ) );
  XNOR2_X1 U1419 ( .A(n880), .B(n879), .ZN(n882) );
  XNOR2_X1 U1420 ( .A(n882), .B(n881), .ZN(n922) );
  XNOR2_X1 U1421 ( .A(n884), .B(n883), .ZN(n886) );
  XNOR2_X1 U1422 ( .A(n886), .B(n885), .ZN(n921) );
  INV_X1 U1423 ( .A(n922), .ZN(n900) );
  NAND2_X1 U1424 ( .A1(n1478), .A2(b[19]), .ZN(n888) );
  NAND2_X1 U1425 ( .A1(n1579), .A2(b[18]), .ZN(n887) );
  OAI211_X1 U1426 ( .C1(b[18]), .C2(n1481), .A(n888), .B(n887), .ZN(n889) );
  AOI21_X1 U1427 ( .B1(n1583), .B2(n1341), .A(n889), .ZN(n994) );
  OAI21_X1 U1428 ( .B1(n1684), .B2(n1694), .A(n994), .ZN(n890) );
  OAI211_X1 U1429 ( .C1(b[9]), .C2(b[8]), .A(n890), .B(a[23]), .ZN(n956) );
  INV_X1 U1430 ( .A(n956), .ZN(n899) );
  NOR2_X1 U1431 ( .A1(n1437), .A2(n1247), .ZN(n892) );
  NOR2_X1 U1432 ( .A1(n1434), .A2(n893), .ZN(n891) );
  AOI211_X1 U1433 ( .C1(n1531), .C2(n893), .A(n892), .B(n891), .ZN(n894) );
  OAI21_X1 U1434 ( .B1(b[18]), .B2(n1394), .A(n894), .ZN(n953) );
  NOR2_X1 U1435 ( .A1(n1449), .A2(b[16]), .ZN(n896) );
  MUX2_X1 U1436 ( .A(n1902), .B(n1439), .S(n1131), .Z(n895) );
  AOI211_X1 U1437 ( .C1(b[16]), .C2(n989), .A(n896), .B(n895), .ZN(n954) );
  OAI21_X1 U1438 ( .B1(n956), .B2(n897), .A(n954), .ZN(n898) );
  OAI21_X1 U1439 ( .B1(n899), .B2(n953), .A(n898), .ZN(n923) );
  OAI21_X1 U1440 ( .B1(n921), .B2(n900), .A(n923), .ZN(n901) );
  OAI21_X1 U1441 ( .B1(n922), .B2(n902), .A(n901), .ZN(\intadd_60/A[2] ) );
  OAI22_X1 U1442 ( .A1(b[21]), .A2(n1596), .B1(n1619), .B2(n1996), .ZN(n904)
         );
  NOR2_X1 U1443 ( .A1(n1616), .A2(b[22]), .ZN(n903) );
  AOI211_X1 U1444 ( .C1(n1617), .C2(b[21]), .A(n904), .B(n903), .ZN(n927) );
  NAND2_X1 U1445 ( .A1(a[23]), .A2(b[10]), .ZN(n925) );
  NOR2_X1 U1446 ( .A1(n927), .A2(n905), .ZN(n908) );
  NAND2_X1 U1447 ( .A1(n1725), .A2(b[23]), .ZN(n906) );
  OAI211_X1 U1448 ( .C1(b[23]), .C2(n1730), .A(n1722), .B(n906), .ZN(n926) );
  OAI22_X1 U1449 ( .A1(n908), .A2(n926), .B1(n907), .B2(n925), .ZN(
        \intadd_60/A[1] ) );
  INV_X1 U1450 ( .A(n909), .ZN(n911) );
  NAND2_X1 U1451 ( .A1(n911), .A2(n910), .ZN(n913) );
  XOR2_X1 U1452 ( .A(n913), .B(n912), .Z(\intadd_60/B[2] ) );
  AOI21_X1 U1453 ( .B1(b[11]), .B2(b[10]), .A(n914), .ZN(n915) );
  XOR2_X1 U1454 ( .A(n916), .B(n915), .Z(\intadd_60/B[1] ) );
  AND2_X1 U1455 ( .A1(n1893), .A2(b[12]), .ZN(n920) );
  NOR2_X1 U1456 ( .A1(n1994), .A2(b[12]), .ZN(n919) );
  NAND2_X1 U1457 ( .A1(n1999), .A2(b[11]), .ZN(n917) );
  OAI21_X1 U1458 ( .B1(n1895), .B2(b[11]), .A(n917), .ZN(n918) );
  NOR3_X1 U1459 ( .A1(n920), .A2(n919), .A3(n918), .ZN(\intadd_60/B[0] ) );
  XNOR2_X1 U1460 ( .A(n922), .B(n921), .ZN(n924) );
  XOR2_X1 U1461 ( .A(n924), .B(n923), .Z(\intadd_59/A[2] ) );
  XOR2_X1 U1462 ( .A(n926), .B(n925), .Z(n928) );
  XOR2_X1 U1463 ( .A(n928), .B(n927), .Z(\intadd_59/A[1] ) );
  MUX2_X1 U1464 ( .A(n1262), .B(n1450), .S(n1602), .Z(n929) );
  OAI21_X1 U1465 ( .B1(n1131), .B2(n1448), .A(n929), .ZN(n930) );
  AOI21_X1 U1466 ( .B1(n1900), .B2(n1131), .A(n930), .ZN(\intadd_59/A[0] ) );
  NOR2_X1 U1467 ( .A1(n1994), .A2(b[11]), .ZN(n932) );
  MUX2_X1 U1468 ( .A(n1999), .B(n1869), .S(n1732), .Z(n931) );
  AOI211_X1 U1469 ( .C1(b[11]), .C2(n1893), .A(n932), .B(n931), .ZN(n943) );
  AOI22_X1 U1470 ( .A1(b[17]), .A2(n1437), .B1(n1394), .B2(n893), .ZN(n933) );
  AOI21_X1 U1471 ( .B1(n1531), .B2(n1246), .A(n933), .ZN(n934) );
  OAI21_X1 U1472 ( .B1(n1434), .B2(n1246), .A(n934), .ZN(n941) );
  INV_X1 U1473 ( .A(n941), .ZN(n935) );
  NOR2_X1 U1474 ( .A1(n943), .A2(n935), .ZN(n937) );
  NAND2_X1 U1475 ( .A1(n1251), .A2(a[9]), .ZN(n940) );
  OAI22_X1 U1476 ( .A1(n937), .A2(n940), .B1(n936), .B2(n941), .ZN(
        \intadd_59/B[1] ) );
  MUX2_X1 U1477 ( .A(n1703), .B(n1702), .S(n1996), .Z(n938) );
  OAI21_X1 U1478 ( .B1(n1723), .B2(n2165), .A(n938), .ZN(n939) );
  AOI21_X1 U1479 ( .B1(n1689), .B2(n2165), .A(n939), .ZN(\intadd_59/B[0] ) );
  XNOR2_X1 U1480 ( .A(n941), .B(n940), .ZN(n942) );
  XNOR2_X1 U1481 ( .A(n943), .B(n942), .ZN(\intadd_48/A[2] ) );
  AND2_X1 U1482 ( .A1(n1531), .A2(n1602), .ZN(n944) );
  AOI21_X1 U1483 ( .B1(b[14]), .B2(n1530), .A(n944), .ZN(n946) );
  NAND2_X1 U1484 ( .A1(n1529), .A2(b[15]), .ZN(n945) );
  OAI211_X1 U1485 ( .C1(b[15]), .C2(n1394), .A(n946), .B(n945), .ZN(n1063) );
  INV_X1 U1486 ( .A(n1063), .ZN(n949) );
  NOR2_X1 U1487 ( .A1(n1994), .A2(b[9]), .ZN(n948) );
  MUX2_X1 U1488 ( .A(n1999), .B(n1869), .S(n1694), .Z(n947) );
  AOI211_X1 U1489 ( .C1(b[9]), .C2(n1893), .A(n948), .B(n947), .ZN(n1064) );
  OAI21_X1 U1490 ( .B1(n1062), .B2(n949), .A(n1064), .ZN(n950) );
  OAI21_X1 U1491 ( .B1(n1063), .B2(n1771), .A(n950), .ZN(\intadd_48/A[1] ) );
  OAI22_X1 U1492 ( .A1(n1596), .A2(b[18]), .B1(n1619), .B2(n1341), .ZN(n952)
         );
  NOR2_X1 U1493 ( .A1(n1616), .A2(b[19]), .ZN(n951) );
  AOI211_X1 U1494 ( .C1(n1617), .C2(b[18]), .A(n952), .B(n951), .ZN(
        \intadd_48/A[0] ) );
  XNOR2_X1 U1495 ( .A(n954), .B(n953), .ZN(n955) );
  XOR2_X1 U1496 ( .A(n956), .B(n955), .Z(n1018) );
  INV_X1 U1497 ( .A(n1018), .ZN(n981) );
  INV_X1 U1498 ( .A(\intadd_60/SUM[0] ), .ZN(n980) );
  NOR2_X1 U1499 ( .A1(n1481), .A2(b[17]), .ZN(n957) );
  AOI21_X1 U1500 ( .B1(n1579), .B2(b[17]), .A(n957), .ZN(n960) );
  NAND2_X1 U1501 ( .A1(n1583), .A2(n1247), .ZN(n959) );
  NAND2_X1 U1502 ( .A1(n1478), .A2(b[18]), .ZN(n958) );
  NAND3_X1 U1503 ( .A1(n960), .A2(n959), .A3(n958), .ZN(n1009) );
  AOI22_X1 U1504 ( .A1(n1389), .A2(b[20]), .B1(n1618), .B2(n1341), .ZN(n962)
         );
  NAND2_X1 U1505 ( .A1(n1617), .A2(b[19]), .ZN(n961) );
  OAI211_X1 U1506 ( .C1(b[20]), .C2(n1616), .A(n962), .B(n961), .ZN(n1010) );
  MUX2_X1 U1507 ( .A(n1999), .B(n1869), .S(n1684), .Z(n963) );
  AOI21_X1 U1508 ( .B1(n1893), .B2(b[10]), .A(n963), .ZN(n964) );
  OAI21_X1 U1509 ( .B1(b[10]), .B2(n1994), .A(n964), .ZN(n1011) );
  FA_X1 U1510 ( .A(n1009), .B(n1010), .CI(n1011), .CO(n1001), .S() );
  NOR2_X1 U1511 ( .A1(n1722), .A2(b[22]), .ZN(n968) );
  NAND2_X1 U1512 ( .A1(n1725), .A2(b[21]), .ZN(n965) );
  OAI21_X1 U1513 ( .B1(n1702), .B2(b[21]), .A(n965), .ZN(n967) );
  NOR2_X1 U1514 ( .A1(n1723), .A2(n1996), .ZN(n966) );
  NOR3_X1 U1515 ( .A1(n968), .A2(n967), .A3(n966), .ZN(n1015) );
  AOI21_X1 U1518 ( .B1(n1742), .B2(b[23]), .A(n970), .ZN(n971) );
  NAND2_X1 U1519 ( .A1(n1698), .A2(n971), .ZN(n1014) );
  NAND2_X1 U1520 ( .A1(a[23]), .A2(b[8]), .ZN(n1013) );
  NAND2_X1 U1521 ( .A1(n1014), .A2(n1013), .ZN(n977) );
  NOR2_X1 U1522 ( .A1(n1616), .A2(b[21]), .ZN(n975) );
  NAND2_X1 U1523 ( .A1(n1617), .A2(b[20]), .ZN(n973) );
  NAND2_X1 U1524 ( .A1(n1618), .A2(n1309), .ZN(n972) );
  OAI211_X1 U1525 ( .C1(n1991), .C2(n1619), .A(n973), .B(n972), .ZN(n974) );
  NOR2_X1 U1526 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1527 ( .A1(n1014), .A2(n1013), .ZN(n978) );
  AOI211_X1 U1528 ( .C1(n1015), .C2(n977), .A(n976), .B(n978), .ZN(n997) );
  OAI211_X1 U1529 ( .C1(n1015), .C2(n978), .A(n977), .B(n976), .ZN(n998) );
  OAI21_X1 U1530 ( .B1(n1001), .B2(n997), .A(n998), .ZN(n1019) );
  OAI21_X1 U1531 ( .B1(\intadd_60/SUM[0] ), .B2(n1018), .A(n1019), .ZN(n979)
         );
  OAI21_X1 U1532 ( .B1(n981), .B2(n980), .A(n979), .ZN(\intadd_48/B[4] ) );
  AOI22_X1 U1533 ( .A1(b[16]), .A2(n1437), .B1(n1394), .B2(n1246), .ZN(n982)
         );
  AOI21_X1 U1534 ( .B1(n1531), .B2(n1131), .A(n982), .ZN(n983) );
  OAI21_X1 U1535 ( .B1(n1434), .B2(n1131), .A(n983), .ZN(n1005) );
  NOR2_X1 U1536 ( .A1(n1883), .A2(n1717), .ZN(n984) );
  AOI21_X1 U1537 ( .B1(n1377), .B2(n1717), .A(n984), .ZN(n987) );
  NAND2_X1 U1538 ( .A1(n1884), .A2(n1273), .ZN(n986) );
  NAND2_X1 U1539 ( .A1(n1374), .A2(b[12]), .ZN(n985) );
  NAND3_X1 U1540 ( .A1(n987), .A2(n986), .A3(n985), .ZN(n1007) );
  MUX2_X1 U1541 ( .A(n1902), .B(n1439), .S(n1670), .Z(n988) );
  AOI21_X1 U1542 ( .B1(n989), .B2(b[14]), .A(n988), .ZN(n990) );
  OAI21_X1 U1543 ( .B1(b[14]), .B2(n1449), .A(n990), .ZN(n1006) );
  FA_X1 U1544 ( .A(n1005), .B(n1007), .CI(n1006), .CO(n1022), .S() );
  INV_X1 U1545 ( .A(\intadd_59/SUM[0] ), .ZN(n996) );
  NOR2_X1 U1546 ( .A1(\intadd_59/SUM[0] ), .A2(n991), .ZN(n995) );
  XOR2_X1 U1549 ( .A(n994), .B(n993), .Z(n1021) );
  OAI22_X1 U1550 ( .A1(n1022), .A2(n996), .B1(n995), .B2(n1021), .ZN(
        \intadd_48/B[3] ) );
  INV_X1 U1551 ( .A(n997), .ZN(n999) );
  NAND2_X1 U1552 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1553 ( .A(n1001), .B(n1000), .Z(\intadd_48/B[2] ) );
  INV_X1 U1554 ( .A(n1030), .ZN(n1069) );
  AOI21_X1 U1555 ( .B1(b[7]), .B2(n1069), .A(n1002), .ZN(\intadd_48/B[1] ) );
  MUX2_X1 U1556 ( .A(n1262), .B(n1450), .S(n1273), .Z(n1003) );
  OAI21_X1 U1557 ( .B1(n1670), .B2(n1448), .A(n1003), .ZN(n1004) );
  AOI21_X1 U1558 ( .B1(n1900), .B2(n1670), .A(n1004), .ZN(\intadd_48/B[0] ) );
  XOR2_X1 U1559 ( .A(n1006), .B(n1005), .Z(n1008) );
  XOR2_X1 U1560 ( .A(n1008), .B(n1007), .Z(n1060) );
  XOR2_X1 U1561 ( .A(n1010), .B(n1009), .Z(n1012) );
  XOR2_X1 U1562 ( .A(n1012), .B(n1011), .Z(n1059) );
  XNOR2_X1 U1563 ( .A(n1014), .B(n1013), .ZN(n1016) );
  XOR2_X1 U1564 ( .A(n1016), .B(n1015), .Z(n1058) );
  AND2_X1 U1565 ( .A1(n1059), .A2(n1058), .ZN(n1017) );
  OAI22_X1 U1566 ( .A1(n1060), .A2(n1017), .B1(n1059), .B2(n1058), .ZN(
        \intadd_47/A[3] ) );
  XOR2_X1 U1567 ( .A(n1019), .B(n1018), .Z(n1020) );
  XOR2_X1 U1568 ( .A(n1020), .B(\intadd_60/SUM[0] ), .Z(\intadd_47/B[4] ) );
  XOR2_X1 U1569 ( .A(n1022), .B(n1021), .Z(n1023) );
  XOR2_X1 U1570 ( .A(\intadd_59/SUM[0] ), .B(n1023), .Z(\intadd_47/B[3] ) );
  NOR2_X1 U1571 ( .A1(a[6]), .A2(n1024), .ZN(n1025) );
  MUX2_X1 U1572 ( .A(n1025), .B(n1711), .S(b[23]), .Z(n1026) );
  NOR2_X1 U1573 ( .A1(n1026), .A2(n1753), .ZN(n1071) );
  NAND2_X1 U1574 ( .A1(n1741), .A2(n1991), .ZN(n1029) );
  XOR2_X1 U1575 ( .A(a[9]), .B(b[22]), .Z(n1033) );
  NAND2_X1 U1576 ( .A1(n1557), .A2(n1033), .ZN(n1028) );
  NAND2_X1 U1577 ( .A1(n1742), .A2(b[21]), .ZN(n1027) );
  NAND3_X1 U1578 ( .A1(n1029), .A2(n1028), .A3(n1027), .ZN(n1070) );
  NAND2_X1 U1579 ( .A1(n1070), .A2(n1030), .ZN(n1032) );
  INV_X1 U1580 ( .A(n1070), .ZN(n1031) );
  AOI22_X1 U1581 ( .A1(n1071), .A2(n1032), .B1(n1031), .B2(n1069), .ZN(n1077)
         );
  MUX2_X1 U1582 ( .A(n1698), .B(n1697), .S(b[23]), .Z(n1035) );
  OAI21_X1 U1583 ( .B1(n1741), .B2(n1742), .A(n1033), .ZN(n1034) );
  NAND2_X1 U1584 ( .A1(n1035), .A2(n1034), .ZN(n1076) );
  INV_X1 U1585 ( .A(n1076), .ZN(n1041) );
  INV_X1 U1586 ( .A(n1077), .ZN(n1040) );
  NOR2_X1 U1587 ( .A1(n1722), .A2(b[21]), .ZN(n1039) );
  NAND2_X1 U1588 ( .A1(n1725), .A2(b[20]), .ZN(n1036) );
  OAI21_X1 U1589 ( .B1(n1702), .B2(b[20]), .A(n1036), .ZN(n1038) );
  NOR2_X1 U1590 ( .A1(n1723), .A2(n1991), .ZN(n1037) );
  NOR3_X1 U1591 ( .A1(n1039), .A2(n1038), .A3(n1037), .ZN(n1075) );
  OAI21_X1 U1592 ( .B1(n1041), .B2(n1040), .A(n1075), .ZN(n1042) );
  OAI21_X1 U1593 ( .B1(n1077), .B2(n1076), .A(n1042), .ZN(\intadd_47/B[2] ) );
  MUX2_X1 U1594 ( .A(n1262), .B(n1450), .S(n1717), .Z(n1043) );
  OAI21_X1 U1595 ( .B1(n1273), .B2(n1448), .A(n1043), .ZN(n1044) );
  AOI21_X1 U1596 ( .B1(n1900), .B2(n1273), .A(n1044), .ZN(n1104) );
  OAI22_X1 U1597 ( .A1(b[17]), .A2(n1596), .B1(n1619), .B2(n1247), .ZN(n1045)
         );
  AOI21_X1 U1598 ( .B1(b[17]), .B2(n1617), .A(n1045), .ZN(n1046) );
  OAI21_X1 U1599 ( .B1(b[18]), .B2(n1616), .A(n1046), .ZN(n1102) );
  INV_X1 U1600 ( .A(n1102), .ZN(n1047) );
  NOR2_X1 U1601 ( .A1(n1104), .A2(n1047), .ZN(n1051) );
  NAND2_X1 U1602 ( .A1(n1528), .A2(n1602), .ZN(n1049) );
  MUX2_X1 U1603 ( .A(n1435), .B(n1434), .S(b[13]), .Z(n1048) );
  OAI211_X1 U1604 ( .C1(n1602), .C2(n1437), .A(n1049), .B(n1048), .ZN(n1103)
         );
  INV_X1 U1605 ( .A(n1104), .ZN(n1050) );
  OAI22_X1 U1606 ( .A1(n1051), .A2(n1103), .B1(n1050), .B2(n1102), .ZN(
        \intadd_47/B[1] ) );
  MUX2_X1 U1607 ( .A(n1703), .B(n1702), .S(n1341), .Z(n1052) );
  OAI21_X1 U1608 ( .B1(n1309), .B2(n1723), .A(n1052), .ZN(n1053) );
  AOI21_X1 U1609 ( .B1(n1689), .B2(n1309), .A(n1053), .ZN(\intadd_47/B[0] ) );
  AND2_X1 U1610 ( .A1(n1893), .A2(b[8]), .ZN(n1057) );
  NOR2_X1 U1611 ( .A1(n1994), .A2(b[8]), .ZN(n1056) );
  NAND2_X1 U1612 ( .A1(n1999), .A2(b[7]), .ZN(n1054) );
  OAI21_X1 U1613 ( .B1(n1895), .B2(b[7]), .A(n1054), .ZN(n1055) );
  NOR3_X1 U1614 ( .A1(n1057), .A2(n1056), .A3(n1055), .ZN(\intadd_47/CI ) );
  XOR2_X1 U1615 ( .A(n1059), .B(n1058), .Z(n1061) );
  XNOR2_X1 U1616 ( .A(n1061), .B(n1060), .ZN(\intadd_49/A[3] ) );
  XNOR2_X1 U1617 ( .A(n1063), .B(n1062), .ZN(n1065) );
  XOR2_X1 U1618 ( .A(n1065), .B(n1064), .Z(\intadd_49/A[2] ) );
  INV_X1 U1619 ( .A(n1066), .ZN(n1067) );
  NOR2_X1 U1620 ( .A1(n1068), .A2(n1067), .ZN(\intadd_49/A[1] ) );
  XOR2_X1 U1621 ( .A(n1070), .B(n1069), .Z(n1072) );
  XNOR2_X1 U1622 ( .A(n1072), .B(n1071), .ZN(\intadd_71/A[1] ) );
  MUX2_X1 U1623 ( .A(n1712), .B(n1711), .S(b[22]), .Z(n1074) );
  NOR2_X1 U1624 ( .A1(n1769), .A2(b[23]), .ZN(n1073) );
  AOI211_X1 U1625 ( .C1(b[23]), .C2(n1715), .A(n1074), .B(n1073), .ZN(
        \intadd_71/A[0] ) );
  XOR2_X1 U1626 ( .A(n1076), .B(n1075), .Z(n1078) );
  XOR2_X1 U1627 ( .A(n1078), .B(n1077), .Z(\intadd_71/B[2] ) );
  INV_X1 U1628 ( .A(n1083), .ZN(n1081) );
  OAI21_X1 U1629 ( .B1(n1081), .B2(n1080), .A(n1079), .ZN(n1082) );
  OAI21_X1 U1630 ( .B1(n1084), .B2(n1083), .A(n1082), .ZN(\intadd_71/B[1] ) );
  MUX2_X1 U1631 ( .A(n1262), .B(n1450), .S(n1732), .Z(n1085) );
  OAI21_X1 U1632 ( .B1(n1448), .B2(n1717), .A(n1085), .ZN(n1086) );
  AOI21_X1 U1633 ( .B1(n1900), .B2(n1717), .A(n1086), .ZN(\intadd_71/CI ) );
  AND2_X1 U1634 ( .A1(n1893), .A2(b[7]), .ZN(n1090) );
  NOR2_X1 U1635 ( .A1(n1994), .A2(b[7]), .ZN(n1089) );
  NAND2_X1 U1636 ( .A1(n1999), .A2(b[6]), .ZN(n1087) );
  OAI21_X1 U1637 ( .B1(n1895), .B2(b[6]), .A(n1087), .ZN(n1088) );
  NOR3_X1 U1638 ( .A1(n1090), .A2(n1089), .A3(n1088), .ZN(\intadd_49/CI ) );
  INV_X1 U1639 ( .A(n1095), .ZN(n1093) );
  OAI21_X1 U1640 ( .B1(n1093), .B2(n1092), .A(n1091), .ZN(n1094) );
  OAI21_X1 U1641 ( .B1(n1095), .B2(n1136), .A(n1094), .ZN(\intadd_50/A[1] ) );
  MUX2_X1 U1642 ( .A(n1262), .B(n1450), .S(n1684), .Z(n1096) );
  OAI21_X1 U1643 ( .B1(n1732), .B2(n1448), .A(n1096), .ZN(n1097) );
  AOI21_X1 U1644 ( .B1(n1900), .B2(n1732), .A(n1097), .ZN(\intadd_50/A[0] ) );
  INV_X1 U1645 ( .A(\intadd_71/SUM[1] ), .ZN(n1101) );
  NOR2_X1 U1646 ( .A1(\intadd_71/SUM[1] ), .A2(\intadd_49/SUM[1] ), .ZN(n1099)
         );
  OAI22_X1 U1647 ( .A1(n1101), .A2(n1100), .B1(n1099), .B2(n1098), .ZN(
        \intadd_50/B[3] ) );
  XOR2_X1 U1648 ( .A(n1103), .B(n1102), .Z(n1105) );
  XOR2_X1 U1649 ( .A(n1105), .B(n1104), .Z(\intadd_50/B[2] ) );
  NOR2_X1 U1650 ( .A1(n1106), .A2(n1107), .ZN(n1111) );
  INV_X1 U1651 ( .A(n1107), .ZN(n1109) );
  OAI22_X1 U1652 ( .A1(n1111), .A2(n1110), .B1(n1109), .B2(n1108), .ZN(
        \intadd_50/B[1] ) );
  MUX2_X1 U1653 ( .A(n1435), .B(n1434), .S(b[11]), .Z(n1112) );
  OAI21_X1 U1654 ( .B1(n1437), .B2(n1273), .A(n1112), .ZN(n1113) );
  AOI21_X1 U1655 ( .B1(n1528), .B2(n1273), .A(n1113), .ZN(\intadd_50/CI ) );
  INV_X1 U1656 ( .A(n1118), .ZN(n1116) );
  OAI21_X1 U1657 ( .B1(n1116), .B2(n1115), .A(n1114), .ZN(n1117) );
  OAI21_X1 U1658 ( .B1(n1119), .B2(n1118), .A(n1117), .ZN(\intadd_63/A[1] ) );
  MUX2_X1 U1659 ( .A(n1435), .B(n1434), .S(b[10]), .Z(n1120) );
  OAI21_X1 U1660 ( .B1(n1437), .B2(n1717), .A(n1120), .ZN(n1121) );
  AOI21_X1 U1661 ( .B1(n1528), .B2(n1717), .A(n1121), .ZN(\intadd_63/A[0] ) );
  XNOR2_X1 U1662 ( .A(n1123), .B(n1122), .ZN(n1124) );
  XNOR2_X1 U1663 ( .A(\intadd_71/SUM[0] ), .B(n1124), .ZN(n1190) );
  INV_X1 U1664 ( .A(n1190), .ZN(n1129) );
  INV_X1 U1665 ( .A(\intadd_50/SUM[1] ), .ZN(n1128) );
  FA_X1 U1666 ( .A(n1126), .B(n1125), .CI(\intadd_50/SUM[0] ), .CO(n1191), 
        .S() );
  OAI21_X1 U1667 ( .B1(\intadd_50/SUM[1] ), .B2(n1190), .A(n1191), .ZN(n1127)
         );
  OAI21_X1 U1668 ( .B1(n1129), .B2(n1128), .A(n1127), .ZN(\intadd_63/B[3] ) );
  AOI22_X1 U1669 ( .A1(b[16]), .A2(n1619), .B1(n1616), .B2(n1246), .ZN(n1130)
         );
  AOI221_X1 U1670 ( .B1(n1617), .B2(b[15]), .C1(n1618), .C2(n1131), .A(n1130), 
        .ZN(n1144) );
  NAND2_X1 U1671 ( .A1(n1478), .A2(b[14]), .ZN(n1133) );
  NAND2_X1 U1672 ( .A1(n1579), .A2(b[13]), .ZN(n1132) );
  OAI211_X1 U1673 ( .C1(b[13]), .C2(n1481), .A(n1133), .B(n1132), .ZN(n1134)
         );
  AOI21_X1 U1674 ( .B1(n1583), .B2(n1602), .A(n1134), .ZN(n1143) );
  OAI21_X1 U1675 ( .B1(a[23]), .B2(b[4]), .A(n1136), .ZN(n1158) );
  OAI22_X1 U1676 ( .A1(n1187), .A2(n1158), .B1(b[5]), .B2(n1994), .ZN(n1139)
         );
  AOI211_X1 U1677 ( .C1(n1893), .C2(b[5]), .A(n1138), .B(n1139), .ZN(n1142) );
  NAND2_X1 U1678 ( .A1(n1139), .A2(n1138), .ZN(n1140) );
  OAI21_X1 U1679 ( .B1(n1142), .B2(n1141), .A(n1140), .ZN(n1155) );
  NOR2_X1 U1680 ( .A1(n1144), .A2(n1143), .ZN(n1153) );
  AOI21_X1 U1681 ( .B1(n1145), .B2(n1155), .A(n1153), .ZN(\intadd_63/B[2] ) );
  AOI21_X1 U1682 ( .B1(n1147), .B2(n1172), .A(n1146), .ZN(\intadd_63/B[1] ) );
  MUX2_X1 U1683 ( .A(n1262), .B(n1450), .S(n1694), .Z(n1148) );
  OAI21_X1 U1684 ( .B1(n1684), .B2(n1448), .A(n1148), .ZN(n1149) );
  AOI21_X1 U1685 ( .B1(n1900), .B2(n1684), .A(n1149), .ZN(\intadd_63/B[0] ) );
  NOR2_X1 U1686 ( .A1(n1666), .A2(n1247), .ZN(n1151) );
  MUX2_X1 U1687 ( .A(n1739), .B(n1738), .S(b[19]), .Z(n1150) );
  AOI211_X1 U1688 ( .C1(n1741), .C2(n1247), .A(n1151), .B(n1150), .ZN(
        \intadd_63/CI ) );
  NOR2_X1 U1689 ( .A1(n1153), .A2(n1152), .ZN(n1154) );
  XNOR2_X1 U1690 ( .A(n1155), .B(n1154), .ZN(\intadd_61/A[2] ) );
  MUX2_X1 U1691 ( .A(n1703), .B(n1702), .S(n1246), .Z(n1156) );
  OAI21_X1 U1692 ( .B1(n893), .B2(n1723), .A(n1156), .ZN(n1157) );
  AOI21_X1 U1693 ( .B1(n1689), .B2(n893), .A(n1157), .ZN(\intadd_61/A[1] ) );
  OAI22_X1 U1694 ( .A1(n1289), .A2(n1158), .B1(n1895), .B2(b[3]), .ZN(n1159)
         );
  AOI21_X1 U1695 ( .B1(n1999), .B2(b[3]), .A(n1159), .ZN(\intadd_61/A[0] ) );
  INV_X1 U1696 ( .A(n1160), .ZN(n1164) );
  NOR2_X1 U1697 ( .A1(\intadd_63/SUM[1] ), .A2(n1160), .ZN(n1162) );
  OAI22_X1 U1698 ( .A1(n1164), .A2(n1163), .B1(n1162), .B2(n1161), .ZN(
        \intadd_61/B[3] ) );
  INV_X1 U1699 ( .A(n1170), .ZN(n1166) );
  OAI21_X1 U1700 ( .B1(n1167), .B2(n1166), .A(n1165), .ZN(n1168) );
  OAI21_X1 U1701 ( .B1(n1170), .B2(n1169), .A(n1168), .ZN(\intadd_61/B[2] ) );
  OAI211_X1 U1702 ( .C1(n1173), .C2(n2165), .A(n1172), .B(n1186), .ZN(n1175)
         );
  OAI211_X1 U1703 ( .C1(n1176), .C2(n2165), .A(n1175), .B(n1174), .ZN(
        \intadd_61/B[1] ) );
  NAND2_X1 U1704 ( .A1(n1183), .A2(n1996), .ZN(n1177) );
  MUX2_X1 U1705 ( .A(n1996), .B(n1177), .S(a[5]), .Z(n1178) );
  NAND3_X1 U1706 ( .A1(n1178), .A2(n1599), .A3(n1789), .ZN(n1182) );
  OAI21_X1 U1707 ( .B1(b[21]), .B2(n1180), .A(n1179), .ZN(n1181) );
  OAI211_X1 U1708 ( .C1(b[21]), .C2(n1183), .A(n1182), .B(n1181), .ZN(
        \intadd_61/CI ) );
  OAI22_X1 U1709 ( .A1(n1596), .A2(b[13]), .B1(n1619), .B2(n1602), .ZN(n1185)
         );
  NOR2_X1 U1710 ( .A1(n1616), .A2(b[14]), .ZN(n1184) );
  AOI211_X1 U1711 ( .C1(n1617), .C2(b[13]), .A(n1185), .B(n1184), .ZN(
        \intadd_51/A[1] ) );
  OAI21_X1 U1712 ( .B1(a[23]), .B2(b[2]), .A(n1186), .ZN(n1290) );
  NOR2_X1 U1713 ( .A1(n1187), .A2(n1290), .ZN(n1188) );
  AOI211_X1 U1714 ( .C1(b[3]), .C2(n1893), .A(n1189), .B(n1188), .ZN(
        \intadd_51/A[0] ) );
  XNOR2_X1 U1715 ( .A(n1191), .B(n1190), .ZN(n1192) );
  XNOR2_X1 U1716 ( .A(n1192), .B(\intadd_50/SUM[1] ), .ZN(\intadd_51/B[4] ) );
  INV_X1 U1717 ( .A(n1194), .ZN(n1198) );
  INV_X1 U1718 ( .A(n1197), .ZN(n1195) );
  OAI21_X1 U1719 ( .B1(n1195), .B2(n1194), .A(n1193), .ZN(n1196) );
  OAI21_X1 U1720 ( .B1(n1198), .B2(n1197), .A(n1196), .ZN(\intadd_51/B[3] ) );
  OAI22_X1 U1721 ( .A1(n1202), .A2(n1201), .B1(n1200), .B2(n1199), .ZN(
        \intadd_51/B[2] ) );
  MUX2_X1 U1722 ( .A(n1850), .B(n1849), .S(b[23]), .Z(n1204) );
  MUX2_X1 U1723 ( .A(n1852), .B(n1851), .S(b[22]), .Z(n1203) );
  NAND2_X1 U1724 ( .A1(n1204), .A2(n1203), .ZN(n1308) );
  NAND2_X1 U1725 ( .A1(a[23]), .A2(b[1]), .ZN(n1306) );
  OAI21_X1 U1726 ( .B1(n1206), .B2(n1205), .A(n1306), .ZN(n1207) );
  OAI21_X1 U1727 ( .B1(a[1]), .B2(n1308), .A(n1207), .ZN(\intadd_51/B[1] ) );
  MUX2_X1 U1728 ( .A(n1861), .B(n1860), .S(n1991), .Z(n1209) );
  MUX2_X1 U1729 ( .A(n39), .B(n1862), .S(b[20]), .Z(n1208) );
  NOR2_X1 U1730 ( .A1(n1209), .A2(n1208), .ZN(\intadd_51/CI ) );
  XNOR2_X1 U1731 ( .A(n1211), .B(n1210), .ZN(n1213) );
  XNOR2_X1 U1732 ( .A(n1213), .B(n1212), .ZN(\intadd_52/A[4] ) );
  OAI21_X1 U1733 ( .B1(n1216), .B2(n1215), .A(n1214), .ZN(n1217) );
  OAI21_X1 U1734 ( .B1(n1219), .B2(n1218), .A(n1217), .ZN(\intadd_70/A[2] ) );
  MUX2_X1 U1735 ( .A(n1850), .B(n1849), .S(b[20]), .Z(n1221) );
  MUX2_X1 U1736 ( .A(n1852), .B(n1851), .S(b[19]), .Z(n1220) );
  NAND2_X1 U1737 ( .A1(n1221), .A2(n1220), .ZN(n1386) );
  NOR2_X1 U1738 ( .A1(n1722), .A2(b[12]), .ZN(n1225) );
  NAND2_X1 U1739 ( .A1(n1725), .A2(b[11]), .ZN(n1222) );
  OAI21_X1 U1740 ( .B1(n1702), .B2(b[11]), .A(n1222), .ZN(n1224) );
  NOR2_X1 U1741 ( .A1(n1723), .A2(n1273), .ZN(n1223) );
  NOR3_X1 U1742 ( .A1(n1225), .A2(n1224), .A3(n1223), .ZN(n1384) );
  INV_X1 U1743 ( .A(n1384), .ZN(n1230) );
  INV_X1 U1744 ( .A(n1386), .ZN(n1228) );
  OAI22_X1 U1745 ( .A1(b[9]), .A2(n1596), .B1(n1619), .B2(n1732), .ZN(n1227)
         );
  NOR2_X1 U1746 ( .A1(n1616), .A2(b[10]), .ZN(n1226) );
  AOI211_X1 U1747 ( .C1(n1617), .C2(b[9]), .A(n1227), .B(n1226), .ZN(n1385) );
  OAI21_X1 U1748 ( .B1(n1228), .B2(n1384), .A(n1385), .ZN(n1229) );
  OAI21_X1 U1749 ( .B1(n1386), .B2(n1230), .A(n1229), .ZN(\intadd_70/A[1] ) );
  NAND2_X1 U1750 ( .A1(n1231), .A2(b[0]), .ZN(\intadd_70/A[0] ) );
  MUX2_X1 U1751 ( .A(n1703), .B(n1702), .S(n1670), .Z(n1233) );
  NAND2_X1 U1752 ( .A1(n1689), .A2(n1602), .ZN(n1232) );
  OAI211_X1 U1753 ( .C1(n1602), .C2(n1723), .A(n1233), .B(n1232), .ZN(n1359)
         );
  NOR2_X1 U1754 ( .A1(n2167), .A2(b[1]), .ZN(n1236) );
  NOR2_X1 U1755 ( .A1(n1234), .A2(b[0]), .ZN(n1235) );
  OAI21_X1 U1756 ( .B1(n1869), .B2(n1236), .A(n1235), .ZN(n1356) );
  XOR2_X1 U1757 ( .A(n1359), .B(n1356), .Z(n1243) );
  INV_X1 U1758 ( .A(n1239), .ZN(n1237) );
  NAND2_X1 U1759 ( .A1(n1237), .A2(n1238), .ZN(n1242) );
  INV_X1 U1760 ( .A(n1238), .ZN(n1240) );
  AOI22_X1 U1761 ( .A1(n1242), .A2(n1241), .B1(n1240), .B2(n1239), .ZN(n1358)
         );
  XOR2_X1 U1762 ( .A(n1243), .B(n1358), .Z(\intadd_70/B[2] ) );
  MUX2_X1 U1763 ( .A(n1752), .B(n1751), .S(b[15]), .Z(n1245) );
  NAND2_X1 U1764 ( .A1(n1753), .A2(n1246), .ZN(n1244) );
  OAI211_X1 U1765 ( .C1(n1246), .C2(n1770), .A(n1245), .B(n1244), .ZN(n1428)
         );
  MUX2_X1 U1766 ( .A(n144), .B(n1788), .S(n1247), .Z(n1249) );
  MUX2_X1 U1767 ( .A(n1789), .B(n1599), .S(b[17]), .Z(n1248) );
  NAND2_X1 U1768 ( .A1(n1249), .A2(n1248), .ZN(n1430) );
  INV_X1 U1769 ( .A(n1430), .ZN(n1258) );
  INV_X1 U1770 ( .A(n1428), .ZN(n1257) );
  NAND2_X1 U1771 ( .A1(n1250), .A2(b[13]), .ZN(n1253) );
  NOR2_X1 U1772 ( .A1(a[9]), .A2(b[14]), .ZN(n1252) );
  MUX2_X1 U1773 ( .A(n1253), .B(n1252), .S(n1251), .Z(n1254) );
  AOI211_X1 U1774 ( .C1(a[9]), .C2(b[14]), .A(n1255), .B(n1254), .ZN(n1256) );
  AOI21_X1 U1775 ( .B1(n1741), .B2(n1670), .A(n1256), .ZN(n1429) );
  OAI21_X1 U1776 ( .B1(n1258), .B2(n1257), .A(n1429), .ZN(n1259) );
  OAI21_X1 U1777 ( .B1(n1428), .B2(n1430), .A(n1259), .ZN(\intadd_70/B[1] ) );
  MUX2_X1 U1778 ( .A(n1884), .B(n1374), .S(b[2]), .Z(n1261) );
  MUX2_X1 U1779 ( .A(n1375), .B(n1377), .S(n2086), .Z(n1260) );
  NOR2_X1 U1780 ( .A1(n1261), .A2(n1260), .ZN(\intadd_70/B[0] ) );
  MUX2_X1 U1781 ( .A(n1262), .B(n1450), .S(n1787), .Z(n1263) );
  OAI21_X1 U1782 ( .B1(n1651), .B2(n1448), .A(n1263), .ZN(n1264) );
  AOI21_X1 U1783 ( .B1(n1900), .B2(n1651), .A(n1264), .ZN(\intadd_70/CI ) );
  NOR2_X1 U1784 ( .A1(n1481), .A2(b[9]), .ZN(n1265) );
  AOI21_X1 U1785 ( .B1(n1579), .B2(b[9]), .A(n1265), .ZN(n1268) );
  NAND2_X1 U1786 ( .A1(n1583), .A2(n1732), .ZN(n1267) );
  NAND2_X1 U1787 ( .A1(n1478), .A2(b[10]), .ZN(n1266) );
  NAND3_X1 U1788 ( .A1(n1268), .A2(n1267), .A3(n1266), .ZN(n1320) );
  INV_X1 U1789 ( .A(n1320), .ZN(n1272) );
  AOI22_X1 U1790 ( .A1(b[16]), .A2(n1697), .B1(n1698), .B2(n1246), .ZN(n1269)
         );
  OAI21_X1 U1791 ( .B1(n1701), .B2(b[15]), .A(n1270), .ZN(n1271) );
  AOI21_X1 U1792 ( .B1(n1742), .B2(b[15]), .A(n1271), .ZN(n1319) );
  NOR2_X1 U1793 ( .A1(n1272), .A2(n1319), .ZN(n1278) );
  AOI22_X1 U1794 ( .A1(b[12]), .A2(n1619), .B1(n1616), .B2(n1273), .ZN(n1274)
         );
  AOI21_X1 U1795 ( .B1(n1618), .B2(n1717), .A(n1274), .ZN(n1275) );
  OAI21_X1 U1796 ( .B1(n1276), .B2(n1717), .A(n1275), .ZN(n1318) );
  OAI22_X1 U1797 ( .A1(n1278), .A2(n1318), .B1(n1320), .B2(n1277), .ZN(
        \intadd_73/A[1] ) );
  MUX2_X1 U1798 ( .A(n1435), .B(n1434), .S(b[7]), .Z(n1279) );
  OAI21_X1 U1799 ( .B1(n1437), .B2(n1694), .A(n1279), .ZN(n1280) );
  AOI21_X1 U1800 ( .B1(n1528), .B2(n1694), .A(n1280), .ZN(\intadd_73/A[0] ) );
  NAND2_X1 U1801 ( .A1(n1439), .A2(n1611), .ZN(n1282) );
  NAND2_X1 U1802 ( .A1(n1902), .A2(b[5]), .ZN(n1281) );
  OAI211_X1 U1803 ( .C1(n1448), .C2(n1859), .A(n1282), .B(n1281), .ZN(n1284)
         );
  NOR2_X1 U1804 ( .A1(n1449), .A2(b[6]), .ZN(n1283) );
  NOR2_X1 U1805 ( .A1(n1284), .A2(n1283), .ZN(n1314) );
  MUX2_X1 U1806 ( .A(n1850), .B(n1849), .S(b[22]), .Z(n1286) );
  MUX2_X1 U1807 ( .A(n1852), .B(n1851), .S(b[21]), .Z(n1285) );
  NAND2_X1 U1808 ( .A1(n1286), .A2(n1285), .ZN(n1316) );
  INV_X1 U1809 ( .A(n1314), .ZN(n1291) );
  MUX2_X1 U1810 ( .A(n1287), .B(n1895), .S(n2086), .Z(n1288) );
  OAI21_X1 U1811 ( .B1(n1290), .B2(n1289), .A(n1288), .ZN(n1315) );
  AOI21_X1 U1812 ( .B1(n1316), .B2(n1291), .A(n1315), .ZN(n1292) );
  AOI21_X1 U1813 ( .B1(n1314), .B2(n1293), .A(n1292), .ZN(n1326) );
  AOI22_X1 U1814 ( .A1(n1389), .A2(b[13]), .B1(n1618), .B2(n1273), .ZN(n1295)
         );
  NAND2_X1 U1815 ( .A1(n1617), .A2(b[12]), .ZN(n1294) );
  OAI211_X1 U1816 ( .C1(b[13]), .C2(n1616), .A(n1295), .B(n1294), .ZN(n1323)
         );
  INV_X1 U1817 ( .A(n1326), .ZN(n1304) );
  INV_X1 U1818 ( .A(n1323), .ZN(n1303) );
  NOR2_X1 U1819 ( .A1(n1883), .A2(n1787), .ZN(n1296) );
  AOI21_X1 U1820 ( .B1(n1377), .B2(n1787), .A(n1296), .ZN(n1299) );
  NAND2_X1 U1821 ( .A1(n1884), .A2(n1651), .ZN(n1298) );
  NAND2_X1 U1822 ( .A1(n1374), .A2(b[4]), .ZN(n1297) );
  NAND3_X1 U1823 ( .A1(n1299), .A2(n1298), .A3(n1297), .ZN(n1364) );
  OAI21_X1 U1824 ( .B1(n2165), .B2(a[0]), .A(a[1]), .ZN(n1362) );
  NOR2_X1 U1825 ( .A1(n1362), .A2(n1300), .ZN(n1302) );
  INV_X1 U1826 ( .A(n1362), .ZN(n1301) );
  OAI22_X1 U1827 ( .A1(n1364), .A2(n1302), .B1(n1361), .B2(n1301), .ZN(n1324)
         );
  OAI21_X1 U1828 ( .B1(n1304), .B2(n1303), .A(n1324), .ZN(n1305) );
  OAI21_X1 U1829 ( .B1(n1326), .B2(n1323), .A(n1305), .ZN(\intadd_73/B[2] ) );
  XOR2_X1 U1830 ( .A(n1306), .B(a[1]), .Z(n1307) );
  XOR2_X1 U1831 ( .A(n1308), .B(n1307), .Z(\intadd_73/B[1] ) );
  MUX2_X1 U1832 ( .A(n1861), .B(n1860), .S(n1309), .Z(n1311) );
  MUX2_X1 U1833 ( .A(n39), .B(n1862), .S(b[19]), .Z(n1310) );
  NOR2_X1 U1834 ( .A1(n1311), .A2(n1310), .ZN(\intadd_73/B[0] ) );
  MUX2_X1 U1835 ( .A(n1712), .B(n1711), .S(b[17]), .Z(n1313) );
  NOR2_X1 U1836 ( .A1(n1769), .A2(b[18]), .ZN(n1312) );
  AOI211_X1 U1837 ( .C1(n1715), .C2(b[18]), .A(n1313), .B(n1312), .ZN(
        \intadd_73/CI ) );
  XOR2_X1 U1838 ( .A(n1315), .B(n1314), .Z(n1317) );
  XOR2_X1 U1839 ( .A(n1317), .B(n1316), .Z(n1347) );
  XNOR2_X1 U1840 ( .A(n1319), .B(n1318), .ZN(n1321) );
  XNOR2_X1 U1841 ( .A(n1321), .B(n1320), .ZN(n1348) );
  XOR2_X1 U1842 ( .A(n1347), .B(n1351), .Z(n1322) );
  XNOR2_X1 U1843 ( .A(\intadd_73/SUM[0] ), .B(n1322), .ZN(\intadd_52/A[2] ) );
  XOR2_X1 U1844 ( .A(n1324), .B(n1323), .Z(n1325) );
  XOR2_X1 U1845 ( .A(n1326), .B(n1325), .Z(\intadd_62/A[2] ) );
  NAND2_X1 U1846 ( .A1(a[3]), .A2(b[21]), .ZN(n1329) );
  NOR2_X1 U1847 ( .A1(n1331), .A2(b[20]), .ZN(n1328) );
  MUX2_X1 U1848 ( .A(n1329), .B(n1328), .S(n1327), .Z(n1333) );
  AOI21_X1 U1849 ( .B1(n1991), .B2(n1331), .A(n1330), .ZN(n1332) );
  AOI22_X1 U1850 ( .A1(n1333), .A2(n1332), .B1(n1765), .B2(b[20]), .ZN(n1370)
         );
  NOR2_X1 U1854 ( .A1(n1370), .A2(n1336), .ZN(n1340) );
  OAI22_X1 U1855 ( .A1(n1596), .A2(b[10]), .B1(n1619), .B2(n1717), .ZN(n1337)
         );
  AOI21_X1 U1856 ( .B1(b[10]), .B2(n1617), .A(n1337), .ZN(n1338) );
  OAI21_X1 U1857 ( .B1(b[11]), .B2(n1616), .A(n1338), .ZN(n1369) );
  OAI22_X1 U1858 ( .A1(n1340), .A2(n1369), .B1(n1339), .B2(n1368), .ZN(
        \intadd_62/A[1] ) );
  MUX2_X1 U1859 ( .A(n1861), .B(n1860), .S(n1341), .Z(n1343) );
  MUX2_X1 U1860 ( .A(n39), .B(n1862), .S(b[18]), .Z(n1342) );
  NOR2_X1 U1861 ( .A1(n1343), .A2(n1342), .ZN(\intadd_62/A[0] ) );
  XOR2_X1 U1862 ( .A(n1345), .B(n1344), .Z(n1346) );
  XOR2_X1 U1863 ( .A(\intadd_51/SUM[0] ), .B(n1346), .Z(n1420) );
  INV_X1 U1864 ( .A(\intadd_73/SUM[0] ), .ZN(n1350) );
  OAI21_X1 U1865 ( .B1(\intadd_73/SUM[0] ), .B2(n1348), .A(n1347), .ZN(n1349)
         );
  OAI21_X1 U1866 ( .B1(n1351), .B2(n1350), .A(n1349), .ZN(n1419) );
  OAI21_X1 U1867 ( .B1(\intadd_73/SUM[1] ), .B2(n1420), .A(n1419), .ZN(n1352)
         );
  OAI21_X1 U1868 ( .B1(n1354), .B2(n1353), .A(n1352), .ZN(\intadd_62/B[3] ) );
  INV_X1 U1869 ( .A(n1358), .ZN(n1355) );
  NOR2_X1 U1870 ( .A1(n1355), .A2(n1356), .ZN(n1360) );
  OAI22_X1 U1871 ( .A1(n1360), .A2(n1359), .B1(n1358), .B2(n1357), .ZN(
        \intadd_62/B[2] ) );
  XNOR2_X1 U1872 ( .A(n1362), .B(n1361), .ZN(n1363) );
  XNOR2_X1 U1873 ( .A(n1364), .B(n1363), .ZN(\intadd_62/B[1] ) );
  MUX2_X1 U1874 ( .A(n1435), .B(n1434), .S(b[6]), .Z(n1365) );
  OAI21_X1 U1875 ( .B1(n1437), .B2(n1735), .A(n1365), .ZN(n1366) );
  AOI21_X1 U1876 ( .B1(n1528), .B2(n1735), .A(n1366), .ZN(\intadd_62/B[0] ) );
  MUX2_X1 U1877 ( .A(n1865), .B(n2083), .S(b[22]), .Z(n1367) );
  AOI21_X1 U1878 ( .B1(n1867), .B2(n1991), .A(n1367), .ZN(\intadd_52/A[0] ) );
  XOR2_X1 U1879 ( .A(n1369), .B(n1368), .Z(n1371) );
  XOR2_X1 U1880 ( .A(n1371), .B(n1370), .Z(\intadd_52/B[1] ) );
  MUX2_X1 U1881 ( .A(n1435), .B(n1434), .S(b[5]), .Z(n1372) );
  OAI21_X1 U1882 ( .B1(n1437), .B2(n1859), .A(n1372), .ZN(n1373) );
  AOI21_X1 U1883 ( .B1(n1528), .B2(n1859), .A(n1373), .ZN(\intadd_52/B[0] ) );
  MUX2_X1 U1884 ( .A(n1884), .B(n1374), .S(b[1]), .Z(n1378) );
  INV_X1 U1885 ( .A(n2009), .ZN(n2012) );
  MUX2_X1 U1886 ( .A(n2012), .B(n1375), .S(b[0]), .Z(n1376) );
  NOR3_X1 U1887 ( .A1(n1378), .A2(n1377), .A3(n1376), .ZN(n1381) );
  NOR2_X1 U1888 ( .A1(n1381), .A2(n1380), .ZN(\intadd_80/A[1] ) );
  MUX2_X1 U1889 ( .A(n1449), .B(n1448), .S(b[2]), .Z(n1383) );
  MUX2_X1 U1890 ( .A(n1262), .B(n1450), .S(n2086), .Z(n1382) );
  NAND2_X1 U1891 ( .A1(n1383), .A2(n1382), .ZN(\intadd_80/A[0] ) );
  XNOR2_X1 U1892 ( .A(n1385), .B(n1384), .ZN(n1387) );
  XNOR2_X1 U1893 ( .A(n1387), .B(n1386), .ZN(\intadd_80/B[2] ) );
  MUX2_X1 U1894 ( .A(n1618), .B(n1617), .S(b[8]), .Z(n1388) );
  AOI21_X1 U1895 ( .B1(n1389), .B2(b[9]), .A(n1388), .ZN(n1390) );
  OAI21_X1 U1896 ( .B1(b[9]), .B2(n1616), .A(n1390), .ZN(\intadd_80/B[1] ) );
  NOR2_X1 U1897 ( .A1(n1391), .A2(n2084), .ZN(\intadd_80/B[0] ) );
  MUX2_X1 U1898 ( .A(n1531), .B(n1530), .S(b[3]), .Z(n1392) );
  AOI21_X1 U1899 ( .B1(b[4]), .B2(n1529), .A(n1392), .ZN(n1393) );
  OAI21_X1 U1900 ( .B1(b[4]), .B2(n1394), .A(n1393), .ZN(\intadd_80/CI ) );
  INV_X1 U1902 ( .A(n1396), .ZN(n1397) );
  NOR2_X1 U1903 ( .A1(n1398), .A2(n1397), .ZN(n1412) );
  AOI211_X1 U1904 ( .C1(n1415), .C2(n1413), .A(n1414), .B(n1412), .ZN(n1571)
         );
  NOR2_X1 U1906 ( .A1(n1701), .A2(b[10]), .ZN(n1399) );
  NOR2_X1 U1908 ( .A1(n1437), .A2(n1787), .ZN(n1402) );
  AOI21_X1 U1909 ( .B1(n1528), .B2(n1787), .A(n1402), .ZN(n1404) );
  MUX2_X1 U1910 ( .A(n1435), .B(n1434), .S(b[2]), .Z(n1403) );
  NAND2_X1 U1911 ( .A1(n1404), .A2(n1403), .ZN(n1575) );
  NOR2_X1 U1912 ( .A1(n1481), .A2(b[4]), .ZN(n1405) );
  AOI21_X1 U1913 ( .B1(n1579), .B2(b[4]), .A(n1405), .ZN(n1408) );
  NAND2_X1 U1914 ( .A1(n1583), .A2(n1611), .ZN(n1407) );
  NAND2_X1 U1915 ( .A1(n1478), .A2(b[5]), .ZN(n1406) );
  NAND3_X1 U1916 ( .A1(n1408), .A2(n1407), .A3(n1406), .ZN(n1409) );
  NAND2_X1 U1917 ( .A1(n1575), .A2(n1409), .ZN(n1411) );
  AOI22_X1 U1918 ( .A1(n1576), .A2(n1411), .B1(n1574), .B2(n1410), .ZN(n1572)
         );
  NOR2_X1 U1919 ( .A1(n1571), .A2(n1572), .ZN(n1418) );
  INV_X1 U1920 ( .A(n1412), .ZN(n1417) );
  OAI21_X1 U1921 ( .B1(n1415), .B2(n1414), .A(n1413), .ZN(n1416) );
  NOR2_X1 U1922 ( .A1(n1417), .A2(n1416), .ZN(n1570) );
  NOR2_X1 U1923 ( .A1(n1418), .A2(n1570), .ZN(\intadd_78/A[1] ) );
  XNOR2_X1 U1924 ( .A(n1420), .B(n1419), .ZN(n1421) );
  XNOR2_X1 U1925 ( .A(\intadd_73/SUM[1] ), .B(n1421), .ZN(\intadd_53/A[4] ) );
  NOR2_X1 U1926 ( .A1(n1422), .A2(n1423), .ZN(n1427) );
  INV_X1 U1927 ( .A(n1422), .ZN(n1425) );
  OAI22_X1 U1928 ( .A1(n1427), .A2(n1426), .B1(n1425), .B2(n1424), .ZN(
        \intadd_53/A[3] ) );
  XOR2_X1 U1929 ( .A(n1429), .B(n1428), .Z(n1431) );
  XOR2_X1 U1930 ( .A(n1431), .B(n1430), .Z(\intadd_53/A[1] ) );
  NOR2_X1 U1931 ( .A1(n1666), .A2(n1273), .ZN(n1433) );
  MUX2_X1 U1932 ( .A(n1739), .B(n1738), .S(b[13]), .Z(n1432) );
  AOI211_X1 U1933 ( .C1(n1741), .C2(n1273), .A(n1433), .B(n1432), .ZN(
        \intadd_53/A[0] ) );
  MUX2_X1 U1934 ( .A(n1435), .B(n1434), .S(b[4]), .Z(n1436) );
  OAI21_X1 U1935 ( .B1(n1611), .B2(n1437), .A(n1436), .ZN(n1438) );
  AOI21_X1 U1936 ( .B1(n1528), .B2(n1611), .A(n1438), .ZN(\intadd_53/B[0] ) );
  NOR2_X1 U1937 ( .A1(n1448), .A2(n1787), .ZN(n1441) );
  MUX2_X1 U1938 ( .A(n1902), .B(n1439), .S(n1740), .Z(n1440) );
  AOI211_X1 U1939 ( .C1(n1900), .C2(n1787), .A(n1441), .B(n1440), .ZN(
        \intadd_53/CI ) );
  XNOR2_X1 U1941 ( .A(n1445), .B(n1444), .ZN(n1447) );
  XNOR2_X1 U1942 ( .A(n1447), .B(n1446), .ZN(n1498) );
  MUX2_X1 U1943 ( .A(n1449), .B(n1448), .S(b[1]), .Z(n1452) );
  MUX2_X1 U1944 ( .A(n1262), .B(n1450), .S(n2084), .Z(n1451) );
  NAND2_X1 U1945 ( .A1(n1452), .A2(n1451), .ZN(n1526) );
  MUX2_X1 U1946 ( .A(n144), .B(n1788), .S(n1246), .Z(n1456) );
  MUX2_X1 U1947 ( .A(n1789), .B(n1599), .S(b[15]), .Z(n1455) );
  NOR2_X1 U1948 ( .A1(n1770), .A2(n1602), .ZN(n1459) );
  NOR2_X1 U1949 ( .A1(n1769), .A2(b[14]), .ZN(n1458) );
  MUX2_X1 U1950 ( .A(n1712), .B(n1711), .S(b[13]), .Z(n1457) );
  NOR3_X1 U1951 ( .A1(n1459), .A2(n1458), .A3(n1457), .ZN(n1460) );
  NAND2_X1 U1952 ( .A1(n1501), .A2(n1460), .ZN(n1462) );
  AOI22_X1 U1953 ( .A1(n1524), .A2(n1462), .B1(n1500), .B2(n1461), .ZN(n1496)
         );
  NOR2_X1 U1954 ( .A1(n1463), .A2(n1496), .ZN(n1469) );
  XOR2_X1 U1955 ( .A(n1465), .B(n1464), .Z(n1467) );
  XNOR2_X1 U1956 ( .A(n1467), .B(n1466), .ZN(n1497) );
  OAI22_X1 U1957 ( .A1(n1469), .A2(n1497), .B1(n1498), .B2(n1468), .ZN(
        \intadd_79/A[2] ) );
  NOR2_X1 U1958 ( .A1(n1666), .A2(n1717), .ZN(n1471) );
  MUX2_X1 U1959 ( .A(n1739), .B(n1738), .S(b[12]), .Z(n1470) );
  AOI211_X1 U1960 ( .C1(n1741), .C2(n1717), .A(n1471), .B(n1470), .ZN(
        \intadd_79/A[0] ) );
  INV_X1 U1961 ( .A(n1472), .ZN(n1474) );
  NAND2_X1 U1962 ( .A1(n1474), .A2(n1473), .ZN(n1476) );
  XOR2_X1 U1963 ( .A(n1476), .B(n1475), .Z(\intadd_79/B[2] ) );
  MUX2_X1 U1964 ( .A(n1856), .B(n1855), .S(b[20]), .Z(n1477) );
  OAI21_X1 U1965 ( .B1(b[19]), .B2(n1858), .A(n1477), .ZN(n1492) );
  NAND2_X1 U1966 ( .A1(n1478), .A2(b[6]), .ZN(n1480) );
  NAND2_X1 U1967 ( .A1(n1579), .A2(b[5]), .ZN(n1479) );
  OAI211_X1 U1968 ( .C1(b[5]), .C2(n1481), .A(n1480), .B(n1479), .ZN(n1482) );
  AOI21_X1 U1969 ( .B1(n1583), .B2(n1859), .A(n1482), .ZN(n1493) );
  INV_X1 U1970 ( .A(n1492), .ZN(n1485) );
  OAI22_X1 U1971 ( .A1(b[7]), .A2(n1596), .B1(n1619), .B2(n1694), .ZN(n1484)
         );
  NOR2_X1 U1972 ( .A1(n1616), .A2(b[8]), .ZN(n1483) );
  AOI211_X1 U1973 ( .C1(n1617), .C2(b[7]), .A(n1484), .B(n1483), .ZN(n1494) );
  OAI21_X1 U1974 ( .B1(n1493), .B2(n1485), .A(n1494), .ZN(n1486) );
  OAI21_X1 U1975 ( .B1(n1492), .B2(n1487), .A(n1486), .ZN(\intadd_79/B[1] ) );
  MUX2_X1 U1976 ( .A(n1703), .B(n1702), .S(n1684), .Z(n1488) );
  OAI21_X1 U1977 ( .B1(n1723), .B2(n1732), .A(n1488), .ZN(n1489) );
  AOI21_X1 U1978 ( .B1(n1689), .B2(n1732), .A(n1489), .ZN(\intadd_79/B[0] ) );
  MUX2_X1 U1979 ( .A(n1764), .B(n1763), .S(b[18]), .Z(n1491) );
  MUX2_X1 U1980 ( .A(n1766), .B(n1765), .S(b[17]), .Z(n1490) );
  NOR2_X1 U1981 ( .A1(n1491), .A2(n1490), .ZN(\intadd_79/CI ) );
  XOR2_X1 U1982 ( .A(n1493), .B(n1492), .Z(n1495) );
  XOR2_X1 U1983 ( .A(n1495), .B(n1494), .Z(\intadd_78/CI ) );
  XNOR2_X1 U1984 ( .A(n1497), .B(n1496), .ZN(n1499) );
  XNOR2_X1 U1985 ( .A(n1499), .B(n1498), .ZN(\intadd_56/A[3] ) );
  XOR2_X1 U1986 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR2_X1 U1987 ( .A(n1502), .B(n1524), .Z(\intadd_56/A[2] ) );
  XOR2_X1 U1989 ( .A(a[9]), .B(b[9]), .Z(n1556) );
  NOR2_X1 U1990 ( .A1(n1684), .A2(a[7]), .ZN(n1503) );
  AOI21_X1 U1991 ( .B1(a[8]), .B2(n1684), .A(n1503), .ZN(n1504) );
  NAND2_X1 U1992 ( .A1(n1556), .A2(n1504), .ZN(n1505) );
  OAI22_X1 U1995 ( .A1(n1772), .A2(n1511), .B1(n1510), .B2(n1509), .ZN(n1590)
         );
  INV_X1 U1996 ( .A(n1590), .ZN(n1512) );
  NOR2_X1 U1997 ( .A1(n1592), .A2(n1512), .ZN(n1516) );
  MUX2_X1 U1998 ( .A(n1850), .B(n1849), .S(b[16]), .Z(n1514) );
  MUX2_X1 U1999 ( .A(n1852), .B(n1851), .S(b[15]), .Z(n1513) );
  NAND2_X1 U2000 ( .A1(n1514), .A2(n1513), .ZN(n1591) );
  OAI22_X1 U2001 ( .A1(n1516), .A2(n1591), .B1(n1515), .B2(n1590), .ZN(
        \intadd_56/A[1] ) );
  NAND2_X1 U2002 ( .A1(n1517), .A2(b[0]), .ZN(\intadd_56/A[0] ) );
  INV_X1 U2003 ( .A(n1522), .ZN(n1520) );
  INV_X1 U2004 ( .A(n1523), .ZN(n1519) );
  OAI21_X1 U2005 ( .B1(n1520), .B2(n1519), .A(n1518), .ZN(n1521) );
  OAI21_X1 U2006 ( .B1(n1523), .B2(n1522), .A(n1521), .ZN(\intadd_56/B[2] ) );
  OAI21_X1 U2007 ( .B1(n1527), .B2(n1526), .A(n1525), .ZN(\intadd_56/B[1] ) );
  MUX2_X1 U2008 ( .A(n1529), .B(n1528), .S(n1740), .Z(n1533) );
  MUX2_X1 U2009 ( .A(n1531), .B(n1530), .S(b[1]), .Z(n1532) );
  NOR2_X1 U2010 ( .A1(n1533), .A2(n1532), .ZN(\intadd_56/CI ) );
  XOR2_X1 U2011 ( .A(n1535), .B(n1534), .Z(n1537) );
  XOR2_X1 U2012 ( .A(n1537), .B(n1536), .Z(\intadd_67/B[2] ) );
  MUX2_X1 U2013 ( .A(n1703), .B(n1702), .S(n1611), .Z(n1539) );
  NAND2_X1 U2014 ( .A1(n1689), .A2(n1859), .ZN(n1538) );
  OAI211_X1 U2015 ( .C1(n1859), .C2(n1723), .A(n1539), .B(n1538), .ZN(n1549)
         );
  MUX2_X1 U2016 ( .A(n1856), .B(n1855), .S(b[16]), .Z(n1540) );
  OAI21_X1 U2017 ( .B1(b[15]), .B2(n1858), .A(n1540), .ZN(n1548) );
  MUX2_X1 U2018 ( .A(n1698), .B(n1697), .S(b[8]), .Z(n1542) );
  NAND2_X1 U2019 ( .A1(n1742), .A2(b[7]), .ZN(n1541) );
  OAI211_X1 U2020 ( .C1(b[7]), .C2(n1701), .A(n1542), .B(n1541), .ZN(n1550) );
  OAI22_X1 U2021 ( .A1(n1543), .A2(n1550), .B1(n1549), .B2(n1548), .ZN(
        \intadd_67/B[1] ) );
  MUX2_X1 U2022 ( .A(n1861), .B(n1860), .S(n1273), .Z(n1545) );
  MUX2_X1 U2023 ( .A(n39), .B(n1862), .S(b[11]), .Z(n1544) );
  NOR2_X1 U2024 ( .A1(n1545), .A2(n1544), .ZN(\intadd_67/B[0] ) );
  MUX2_X1 U2025 ( .A(n1712), .B(n1711), .S(b[9]), .Z(n1547) );
  NOR2_X1 U2026 ( .A1(n1769), .A2(b[10]), .ZN(n1546) );
  AOI211_X1 U2027 ( .C1(b[10]), .C2(n1715), .A(n1547), .B(n1546), .ZN(
        \intadd_67/CI ) );
  XOR2_X1 U2028 ( .A(n1549), .B(n1548), .Z(n1551) );
  XOR2_X1 U2029 ( .A(n1551), .B(n1550), .Z(\intadd_76/A[0] ) );
  MUX2_X1 U2030 ( .A(n144), .B(n1788), .S(n1602), .Z(n1553) );
  MUX2_X1 U2031 ( .A(n1789), .B(n1599), .S(b[13]), .Z(n1552) );
  NAND2_X1 U2032 ( .A1(n1553), .A2(n1552), .ZN(n1586) );
  XOR2_X1 U2033 ( .A(n1585), .B(n1586), .Z(n1565) );
  NAND2_X1 U2034 ( .A1(n1742), .A2(b[8]), .ZN(n1554) );
  OAI21_X1 U2035 ( .B1(b[8]), .B2(n1701), .A(n1554), .ZN(n1555) );
  AOI21_X1 U2036 ( .B1(n1557), .B2(n1556), .A(n1555), .ZN(n1567) );
  MUX2_X1 U2037 ( .A(n1850), .B(n1849), .S(b[15]), .Z(n1559) );
  MUX2_X1 U2038 ( .A(n1852), .B(n1851), .S(b[14]), .Z(n1558) );
  NAND2_X1 U2039 ( .A1(n1559), .A2(n1558), .ZN(n1562) );
  NAND2_X1 U2043 ( .A1(n1562), .A2(n1566), .ZN(n1564) );
  INV_X1 U2044 ( .A(n1566), .ZN(n1563) );
  AOI22_X1 U2045 ( .A1(n1567), .A2(n1564), .B1(n1568), .B2(n1563), .ZN(n1589)
         );
  XOR2_X1 U2046 ( .A(n1565), .B(n1589), .Z(\intadd_77/A[1] ) );
  XNOR2_X1 U2047 ( .A(n1567), .B(n1566), .ZN(n1569) );
  XOR2_X1 U2048 ( .A(n1569), .B(n1568), .Z(\intadd_77/A[0] ) );
  NOR2_X1 U2049 ( .A1(n1571), .A2(n1570), .ZN(n1573) );
  XNOR2_X1 U2050 ( .A(n1573), .B(n1572), .ZN(\intadd_55/A[3] ) );
  XOR2_X1 U2051 ( .A(n1575), .B(n1574), .Z(n1577) );
  XNOR2_X1 U2052 ( .A(n1577), .B(n1576), .ZN(\intadd_55/A[2] ) );
  MUX2_X1 U2054 ( .A(n1580), .B(n1579), .S(b[2]), .Z(n1581) );
  AOI211_X1 U2055 ( .C1(n1583), .C2(n1787), .A(n1582), .B(n1581), .ZN(
        \intadd_55/A[0] ) );
  NOR2_X1 U2056 ( .A1(n1585), .A2(n1584), .ZN(n1588) );
  OAI22_X1 U2057 ( .A1(n1589), .A2(n1588), .B1(n1587), .B2(n1586), .ZN(
        \intadd_55/B[2] ) );
  XOR2_X1 U2058 ( .A(n1591), .B(n1590), .Z(n1593) );
  XOR2_X1 U2059 ( .A(n1593), .B(n1592), .Z(\intadd_55/B[1] ) );
  MUX2_X1 U2060 ( .A(n1703), .B(n1702), .S(n1859), .Z(n1594) );
  OAI21_X1 U2061 ( .B1(n1723), .B2(n1735), .A(n1594), .ZN(n1595) );
  AOI21_X1 U2062 ( .B1(n1689), .B2(n1735), .A(n1595), .ZN(\intadd_55/B[0] ) );
  OAI22_X1 U2063 ( .A1(n1596), .A2(b[4]), .B1(n1619), .B2(n1611), .ZN(n1598)
         );
  NOR2_X1 U2064 ( .A1(n1616), .A2(b[5]), .ZN(n1597) );
  AOI211_X1 U2065 ( .C1(n1617), .C2(b[4]), .A(n1598), .B(n1597), .ZN(
        \intadd_55/CI ) );
  MUX2_X1 U2066 ( .A(n144), .B(n1788), .S(n1717), .Z(n1601) );
  MUX2_X1 U2067 ( .A(n1789), .B(n1599), .S(b[10]), .Z(n1600) );
  NAND2_X1 U2068 ( .A1(n1601), .A2(n1600), .ZN(n1663) );
  MUX2_X1 U2072 ( .A(n1698), .B(n1697), .S(b[7]), .Z(n1606) );
  NAND2_X1 U2073 ( .A1(n1742), .A2(b[6]), .ZN(n1605) );
  OAI211_X1 U2074 ( .C1(b[6]), .C2(n1701), .A(n1606), .B(n1605), .ZN(n1664) );
  FA_X1 U2075 ( .A(n1663), .B(n1662), .CI(n1664), .CO(n1661), .S() );
  NOR2_X1 U2076 ( .A1(n1769), .A2(b[9]), .ZN(n1607) );
  AOI21_X1 U2077 ( .B1(b[9]), .B2(n1715), .A(n1607), .ZN(n1609) );
  MUX2_X1 U2078 ( .A(n1752), .B(n1751), .S(b[8]), .Z(n1608) );
  NAND2_X1 U2079 ( .A1(n1609), .A2(n1608), .ZN(n1653) );
  NAND2_X1 U2081 ( .A1(n1725), .A2(b[4]), .ZN(n1610) );
  OAI21_X1 U2082 ( .B1(n1702), .B2(b[4]), .A(n1610), .ZN(n1613) );
  NOR2_X1 U2083 ( .A1(n1723), .A2(n1611), .ZN(n1612) );
  NOR2_X1 U2086 ( .A1(n1653), .A2(n1652), .ZN(n1625) );
  NOR2_X1 U2087 ( .A1(n1616), .A2(b[3]), .ZN(n1622) );
  MUX2_X1 U2088 ( .A(n1618), .B(n1617), .S(b[2]), .Z(n1621) );
  NOR2_X1 U2089 ( .A1(n1619), .A2(n1787), .ZN(n1620) );
  NOR3_X1 U2090 ( .A1(n1622), .A2(n1621), .A3(n1620), .ZN(n1654) );
  INV_X1 U2091 ( .A(n1653), .ZN(n1624) );
  OAI22_X1 U2093 ( .A1(n1625), .A2(n1654), .B1(n1624), .B2(n1623), .ZN(n1628)
         );
  NAND2_X1 U2094 ( .A1(n1628), .A2(n1627), .ZN(n1659) );
  OAI21_X1 U2096 ( .B1(n1661), .B2(n1631), .A(n1658), .ZN(\intadd_77/B[0] ) );
  XNOR2_X1 U2097 ( .A(n1633), .B(n1632), .ZN(n1634) );
  XOR2_X1 U2098 ( .A(n1635), .B(n1634), .Z(\intadd_76/B[1] ) );
  XOR2_X1 U2099 ( .A(n1637), .B(n1636), .Z(n1639) );
  XOR2_X1 U2100 ( .A(n1639), .B(n1638), .Z(\intadd_76/B[0] ) );
  MUX2_X1 U2101 ( .A(n1850), .B(n1849), .S(b[12]), .Z(n1641) );
  MUX2_X1 U2102 ( .A(n1852), .B(n1851), .S(b[11]), .Z(n1640) );
  NAND2_X1 U2103 ( .A1(n1641), .A2(n1640), .ZN(n1691) );
  MUX2_X1 U2104 ( .A(n144), .B(n1788), .S(n1732), .Z(n1643) );
  MUX2_X1 U2105 ( .A(n1789), .B(n1599), .S(b[9]), .Z(n1642) );
  NAND2_X1 U2106 ( .A1(n1643), .A2(n1642), .ZN(n1690) );
  OAI22_X1 U2107 ( .A1(n1644), .A2(n1692), .B1(n1691), .B2(n1690), .ZN(
        \intadd_66/A[2] ) );
  XNOR2_X1 U2108 ( .A(n1646), .B(n1645), .ZN(n1648) );
  XNOR2_X1 U2109 ( .A(n1648), .B(n1647), .ZN(\intadd_66/A[1] ) );
  NOR2_X1 U2110 ( .A1(n1666), .A2(n1651), .ZN(n1650) );
  MUX2_X1 U2111 ( .A(n1739), .B(n1738), .S(b[5]), .Z(n1649) );
  AOI211_X1 U2112 ( .C1(n1741), .C2(n1651), .A(n1650), .B(n1649), .ZN(
        \intadd_66/A[0] ) );
  XNOR2_X1 U2113 ( .A(n1653), .B(n1652), .ZN(n1655) );
  XNOR2_X1 U2114 ( .A(n1655), .B(n1654), .ZN(\intadd_65/A[1] ) );
  MUX2_X1 U2115 ( .A(n1712), .B(n1711), .S(b[7]), .Z(n1657) );
  NOR2_X1 U2116 ( .A1(n1769), .A2(b[8]), .ZN(n1656) );
  AOI211_X1 U2117 ( .C1(b[8]), .C2(n1715), .A(n1657), .B(n1656), .ZN(
        \intadd_65/A[0] ) );
  NAND2_X1 U2118 ( .A1(n1659), .A2(n1658), .ZN(n1660) );
  XOR2_X1 U2119 ( .A(n1661), .B(n1660), .Z(\intadd_65/B[2] ) );
  XNOR2_X1 U2120 ( .A(n1663), .B(n1662), .ZN(n1665) );
  XOR2_X1 U2121 ( .A(n1665), .B(n1664), .Z(\intadd_65/B[1] ) );
  NOR2_X1 U2122 ( .A1(n1666), .A2(n1611), .ZN(n1668) );
  MUX2_X1 U2123 ( .A(n1739), .B(n1738), .S(b[6]), .Z(n1667) );
  AOI211_X1 U2124 ( .C1(n1741), .C2(n1611), .A(n1668), .B(n1667), .ZN(
        \intadd_65/B[0] ) );
  MUX2_X1 U2125 ( .A(n1865), .B(n2083), .S(b[14]), .Z(n1669) );
  AOI21_X1 U2126 ( .B1(n1867), .B2(n1670), .A(n1669), .ZN(\intadd_65/CI ) );
  XOR2_X1 U2127 ( .A(n1672), .B(n1671), .Z(n1673) );
  XNOR2_X1 U2128 ( .A(n1674), .B(n1673), .ZN(\intadd_66/B[2] ) );
  MUX2_X1 U2129 ( .A(n1856), .B(n1855), .S(b[13]), .Z(n1675) );
  OAI21_X1 U2130 ( .B1(b[12]), .B2(n1858), .A(n1675), .ZN(n1718) );
  MUX2_X1 U2131 ( .A(n1850), .B(n1849), .S(b[11]), .Z(n1677) );
  MUX2_X1 U2132 ( .A(n1852), .B(n1851), .S(b[10]), .Z(n1676) );
  NAND2_X1 U2133 ( .A1(n1677), .A2(n1676), .ZN(n1720) );
  INV_X1 U2134 ( .A(n1720), .ZN(n1682) );
  NOR2_X1 U2135 ( .A1(n1770), .A2(n1735), .ZN(n1680) );
  NOR2_X1 U2136 ( .A1(n1769), .A2(b[7]), .ZN(n1679) );
  MUX2_X1 U2137 ( .A(n1712), .B(n1711), .S(b[6]), .Z(n1678) );
  NOR3_X1 U2138 ( .A1(n1680), .A2(n1679), .A3(n1678), .ZN(n1719) );
  OAI21_X1 U2139 ( .B1(n1682), .B2(n1681), .A(n1719), .ZN(n1683) );
  OAI21_X1 U2140 ( .B1(n1718), .B2(n1720), .A(n1683), .ZN(\intadd_66/B[1] ) );
  MUX2_X1 U2141 ( .A(n1861), .B(n1860), .S(n1684), .Z(n1686) );
  MUX2_X1 U2142 ( .A(n39), .B(n1862), .S(b[8]), .Z(n1685) );
  NOR2_X1 U2143 ( .A1(n1686), .A2(n1685), .ZN(\intadd_66/B[0] ) );
  NOR2_X1 U2144 ( .A1(n1723), .A2(n1787), .ZN(n1688) );
  MUX2_X1 U2145 ( .A(n1725), .B(n1726), .S(n1740), .Z(n1687) );
  AOI211_X1 U2146 ( .C1(n1689), .C2(n1787), .A(n1688), .B(n1687), .ZN(
        \intadd_66/CI ) );
  XNOR2_X1 U2147 ( .A(n1691), .B(n1690), .ZN(n1693) );
  XOR2_X1 U2148 ( .A(n1693), .B(n1692), .Z(\intadd_75/A[2] ) );
  MUX2_X1 U2149 ( .A(n1861), .B(n1860), .S(n1694), .Z(n1696) );
  MUX2_X1 U2150 ( .A(n39), .B(n1862), .S(b[7]), .Z(n1695) );
  NOR2_X1 U2151 ( .A1(n1696), .A2(n1695), .ZN(\intadd_75/A[0] ) );
  MUX2_X1 U2152 ( .A(n1698), .B(n1697), .S(b[4]), .Z(n1700) );
  NAND2_X1 U2153 ( .A1(n1742), .A2(b[3]), .ZN(n1699) );
  OAI211_X1 U2154 ( .C1(b[3]), .C2(n1701), .A(n1700), .B(n1699), .ZN(n1746) );
  MUX2_X1 U2155 ( .A(n1723), .B(n1722), .S(n1740), .Z(n1705) );
  MUX2_X1 U2156 ( .A(n1703), .B(n1702), .S(n2086), .Z(n1704) );
  NAND2_X1 U2157 ( .A1(n1705), .A2(n1704), .ZN(n1747) );
  INV_X1 U2158 ( .A(n1747), .ZN(n1708) );
  NAND2_X1 U2159 ( .A1(n1707), .A2(n1706), .ZN(n1745) );
  NOR2_X1 U2160 ( .A1(n1708), .A2(n1745), .ZN(n1710) );
  OAI22_X1 U2161 ( .A1(n1746), .A2(n1710), .B1(n1709), .B2(n1747), .ZN(
        \intadd_75/B[1] ) );
  MUX2_X1 U2162 ( .A(n1712), .B(n1711), .S(b[5]), .Z(n1714) );
  NOR2_X1 U2163 ( .A1(n1769), .A2(b[6]), .ZN(n1713) );
  AOI211_X1 U2164 ( .C1(b[6]), .C2(n1715), .A(n1714), .B(n1713), .ZN(
        \intadd_75/B[0] ) );
  MUX2_X1 U2165 ( .A(n1865), .B(n2083), .S(b[12]), .Z(n1716) );
  AOI21_X1 U2166 ( .B1(n1867), .B2(n1717), .A(n1716), .ZN(\intadd_75/CI ) );
  XNOR2_X1 U2167 ( .A(n1719), .B(n1718), .ZN(n1721) );
  XNOR2_X1 U2168 ( .A(n1721), .B(n1720), .ZN(\intadd_64/A[2] ) );
  MUX2_X1 U2169 ( .A(n1723), .B(n1722), .S(n2086), .Z(n1728) );
  XOR2_X1 U2170 ( .A(a[11]), .B(b[0]), .Z(n1724) );
  OAI21_X1 U2171 ( .B1(n1726), .B2(n1725), .A(n1724), .ZN(n1727) );
  NAND2_X1 U2172 ( .A1(n1728), .A2(n1727), .ZN(n1750) );
  NOR2_X1 U2173 ( .A1(n1730), .A2(n1729), .ZN(n1749) );
  NAND2_X1 U2174 ( .A1(n1750), .A2(n1749), .ZN(\intadd_64/A[1] ) );
  MUX2_X1 U2175 ( .A(n1865), .B(n2083), .S(b[11]), .Z(n1731) );
  AOI21_X1 U2176 ( .B1(n1867), .B2(n1732), .A(n1731), .ZN(\intadd_64/A[0] ) );
  MUX2_X1 U2177 ( .A(n1764), .B(n1763), .S(b[10]), .Z(n1734) );
  MUX2_X1 U2178 ( .A(n1766), .B(n1765), .S(b[9]), .Z(n1733) );
  NOR2_X1 U2179 ( .A1(n1734), .A2(n1733), .ZN(\intadd_64/B[1] ) );
  MUX2_X1 U2180 ( .A(n1861), .B(n1860), .S(n1735), .Z(n1737) );
  MUX2_X1 U2181 ( .A(n39), .B(n1862), .S(b[6]), .Z(n1736) );
  NOR2_X1 U2182 ( .A1(n1737), .A2(n1736), .ZN(\intadd_64/B[0] ) );
  MUX2_X1 U2183 ( .A(n1739), .B(n1738), .S(b[3]), .Z(n1744) );
  MUX2_X1 U2184 ( .A(n1742), .B(n1741), .S(n1740), .Z(n1743) );
  NOR2_X1 U2185 ( .A1(n1744), .A2(n1743), .ZN(\intadd_64/CI ) );
  XNOR2_X1 U2186 ( .A(n1746), .B(n1745), .ZN(n1748) );
  XOR2_X1 U2187 ( .A(n1748), .B(n1747), .Z(\intadd_74/A[1] ) );
  XOR2_X1 U2188 ( .A(n1750), .B(n1749), .Z(\intadd_74/A[0] ) );
  MUX2_X1 U2189 ( .A(n1752), .B(n1751), .S(b[4]), .Z(n1755) );
  NAND2_X1 U2190 ( .A1(n1753), .A2(n1611), .ZN(n1754) );
  OAI211_X1 U2191 ( .C1(n1770), .C2(n1611), .A(n1755), .B(n1754), .ZN(
        \intadd_74/B[0] ) );
  MUX2_X1 U2192 ( .A(n1850), .B(n1849), .S(b[9]), .Z(n1757) );
  MUX2_X1 U2193 ( .A(n1852), .B(n1851), .S(b[8]), .Z(n1756) );
  NAND2_X1 U2194 ( .A1(n1757), .A2(n1756), .ZN(\intadd_74/CI ) );
  INV_X1 U2195 ( .A(n1758), .ZN(n1761) );
  OAI22_X1 U2196 ( .A1(n1762), .A2(n1761), .B1(n1760), .B2(n1759), .ZN(
        \intadd_46/A[1] ) );
  MUX2_X1 U2197 ( .A(n1764), .B(n1763), .S(b[8]), .Z(n1768) );
  MUX2_X1 U2198 ( .A(n1766), .B(n1765), .S(b[7]), .Z(n1767) );
  NOR2_X1 U2199 ( .A1(n1768), .A2(n1767), .ZN(\intadd_46/A[0] ) );
  OAI21_X1 U2200 ( .B1(n1770), .B2(n2086), .A(n1769), .ZN(n1775) );
  MUX2_X1 U2201 ( .A(n1771), .B(n1770), .S(b[1]), .Z(n1773) );
  NAND2_X1 U2202 ( .A1(n1773), .A2(n1772), .ZN(n1774) );
  AOI21_X1 U2205 ( .B1(n1780), .B2(n1779), .A(n1778), .ZN(n1782) );
  NOR2_X1 U2206 ( .A1(n1780), .A2(n1779), .ZN(n1781) );
  NOR2_X1 U2207 ( .A1(n1782), .A2(n1781), .ZN(n1815) );
  XNOR2_X1 U2208 ( .A(n1816), .B(n1815), .ZN(n1793) );
  MUX2_X1 U2209 ( .A(n1850), .B(n1849), .S(b[5]), .Z(n1784) );
  MUX2_X1 U2210 ( .A(n1852), .B(n1851), .S(b[4]), .Z(n1783) );
  MUX2_X1 U2212 ( .A(n1856), .B(n1855), .S(b[7]), .Z(n1786) );
  NAND2_X1 U2213 ( .A1(n1867), .A2(n1859), .ZN(n1785) );
  XNOR2_X1 U2215 ( .A(n1810), .B(n1811), .ZN(n1792) );
  MUX2_X1 U2216 ( .A(n144), .B(n1788), .S(n1787), .Z(n1791) );
  MUX2_X1 U2217 ( .A(n1789), .B(n1599), .S(b[2]), .Z(n1790) );
  NAND2_X1 U2218 ( .A1(n1791), .A2(n1790), .ZN(n1812) );
  XOR2_X1 U2219 ( .A(n1792), .B(n1812), .Z(n1823) );
  XOR2_X1 U2220 ( .A(n1793), .B(n1823), .Z(\intadd_72/A[2] ) );
  MUX2_X1 U2221 ( .A(n1856), .B(n1855), .S(b[5]), .Z(n1794) );
  OAI21_X1 U2222 ( .B1(b[4]), .B2(n1858), .A(n1794), .ZN(\intadd_72/A[0] ) );
  INV_X1 U2223 ( .A(n1797), .ZN(n1795) );
  NOR2_X1 U2224 ( .A1(n1795), .A2(n1796), .ZN(n1800) );
  INV_X1 U2225 ( .A(n1796), .ZN(n1798) );
  OAI22_X1 U2226 ( .A1(n1800), .A2(n1799), .B1(n1798), .B2(n1797), .ZN(
        \intadd_72/B[2] ) );
  MUX2_X1 U2227 ( .A(n1850), .B(n1849), .S(b[3]), .Z(n1803) );
  NAND2_X1 U2228 ( .A1(n1852), .A2(n1740), .ZN(n1801) );
  OAI21_X1 U2229 ( .B1(n1765), .B2(n1740), .A(n1801), .ZN(n1802) );
  NAND2_X1 U2230 ( .A1(n1803), .A2(n1802), .ZN(\intadd_72/CI ) );
  NOR2_X1 U2231 ( .A1(n1816), .A2(n1815), .ZN(n1821) );
  XOR2_X1 U2232 ( .A(n1805), .B(n1804), .Z(n1807) );
  XOR2_X1 U2233 ( .A(n1807), .B(n1806), .Z(n1828) );
  NOR2_X1 U2234 ( .A1(n1809), .A2(n1808), .ZN(n1813) );
  OAI22_X1 U2235 ( .A1(n1813), .A2(n1812), .B1(n1811), .B2(n1810), .ZN(n1827)
         );
  XNOR2_X1 U2236 ( .A(n1828), .B(n1827), .ZN(n1814) );
  XOR2_X1 U2237 ( .A(\intadd_54/SUM[0] ), .B(n1814), .Z(n1820) );
  NAND2_X1 U2238 ( .A1(n1816), .A2(n1815), .ZN(n1822) );
  OAI211_X1 U2239 ( .C1(n1823), .C2(n1821), .A(n1820), .B(n1822), .ZN(n1975)
         );
  NAND2_X1 U2240 ( .A1(\intadd_72/n1 ), .A2(n1975), .ZN(n2052) );
  NOR2_X1 U2241 ( .A1(n1828), .A2(n1827), .ZN(n1817) );
  NOR2_X1 U2242 ( .A1(\intadd_54/SUM[1] ), .A2(n1817), .ZN(n1826) );
  NAND2_X1 U2243 ( .A1(n1828), .A2(n1827), .ZN(n1818) );
  NAND2_X1 U2244 ( .A1(\intadd_54/SUM[0] ), .A2(n1818), .ZN(n1819) );
  NAND2_X1 U2245 ( .A1(n1826), .A2(n1819), .ZN(n2053) );
  INV_X1 U2246 ( .A(n1820), .ZN(n1825) );
  AOI21_X1 U2247 ( .B1(n1823), .B2(n1822), .A(n1821), .ZN(n1824) );
  NAND2_X1 U2248 ( .A1(n1825), .A2(n1824), .ZN(n2051) );
  INV_X1 U2249 ( .A(\intadd_54/SUM[0] ), .ZN(n1829) );
  OAI21_X1 U2250 ( .B1(n1829), .B2(n1828), .A(n1827), .ZN(n1830) );
  OAI211_X1 U2251 ( .C1(n1831), .C2(\intadd_54/SUM[0] ), .A(\intadd_54/SUM[1] ), .B(n1830), .ZN(n2054) );
  OAI211_X1 U2252 ( .C1(n2052), .C2(n1833), .A(n1832), .B(n2054), .ZN(
        \intadd_54/A[2] ) );
  XNOR2_X1 U2253 ( .A(n1835), .B(n1834), .ZN(n1837) );
  XOR2_X1 U2254 ( .A(n1837), .B(n1836), .Z(\intadd_54/A[1] ) );
  INV_X1 U2255 ( .A(\intadd_74/SUM[0] ), .ZN(n1841) );
  OAI21_X1 U2256 ( .B1(n1839), .B2(\intadd_74/SUM[0] ), .A(n1838), .ZN(n1840)
         );
  OAI21_X1 U2257 ( .B1(\intadd_46/SUM[1] ), .B2(n1841), .A(n1840), .ZN(
        \intadd_54/B[4] ) );
  XOR2_X1 U2258 ( .A(\intadd_46/SUM[0] ), .B(n1842), .Z(n1844) );
  XOR2_X1 U2259 ( .A(n1844), .B(n1843), .Z(\intadd_54/B[2] ) );
  XOR2_X1 U2260 ( .A(n1846), .B(n1845), .Z(n1848) );
  XOR2_X1 U2261 ( .A(n1848), .B(n1847), .Z(\intadd_54/B[1] ) );
  MUX2_X1 U2262 ( .A(n1850), .B(n1849), .S(b[6]), .Z(n1854) );
  MUX2_X1 U2263 ( .A(n1852), .B(n1851), .S(b[5]), .Z(n1853) );
  NAND2_X1 U2264 ( .A1(n1854), .A2(n1853), .ZN(\intadd_54/B[0] ) );
  MUX2_X1 U2265 ( .A(n1856), .B(n1855), .S(b[8]), .Z(n1857) );
  OAI21_X1 U2266 ( .B1(b[7]), .B2(n1858), .A(n1857), .ZN(\intadd_54/CI ) );
  MUX2_X1 U2267 ( .A(n1861), .B(n1860), .S(n1859), .Z(n1864) );
  MUX2_X1 U2268 ( .A(n39), .B(n1862), .S(b[5]), .Z(n1863) );
  NOR2_X1 U2269 ( .A1(n1864), .A2(n1863), .ZN(\intadd_46/B[0] ) );
  MUX2_X1 U2270 ( .A(n1865), .B(n2083), .S(b[10]), .Z(n1866) );
  AOI21_X1 U2271 ( .B1(n1867), .B2(n1684), .A(n1866), .ZN(\intadd_46/CI ) );
  XOR2_X1 U2272 ( .A(\intadd_65/SUM[3] ), .B(\intadd_66/n1 ), .Z(n1868) );
  XNOR2_X1 U2273 ( .A(n1907), .B(n1868), .ZN(\d[17]_BAR ) );
  NAND2_X1 U2274 ( .A1(n1869), .A2(n1996), .ZN(n1870) );
  OAI21_X1 U2275 ( .B1(n1994), .B2(b[23]), .A(n1870), .ZN(n1995) );
  INV_X1 U2276 ( .A(n1995), .ZN(n1872) );
  AOI22_X1 U2277 ( .A1(n1893), .A2(b[23]), .B1(n1999), .B2(b[22]), .ZN(n1871)
         );
  NAND2_X1 U2278 ( .A1(n1872), .A2(n1871), .ZN(n1875) );
  NAND2_X1 U2279 ( .A1(a[23]), .A2(b[20]), .ZN(n1992) );
  NAND2_X1 U2280 ( .A1(n1992), .A2(n1991), .ZN(n1998) );
  OAI21_X1 U2281 ( .B1(n2167), .B2(b[20]), .A(b[21]), .ZN(n1873) );
  NAND2_X1 U2282 ( .A1(n1998), .A2(n1873), .ZN(n1874) );
  XOR2_X1 U2283 ( .A(n1875), .B(n1874), .Z(n2013) );
  XOR2_X1 U2284 ( .A(n2013), .B(n2012), .Z(n1889) );
  NAND2_X1 U2285 ( .A1(n1876), .A2(n1996), .ZN(n1880) );
  NAND2_X1 U2286 ( .A1(n1893), .A2(b[22]), .ZN(n1879) );
  NOR2_X1 U2287 ( .A1(n1895), .A2(b[21]), .ZN(n1877) );
  AOI21_X1 U2288 ( .B1(n1999), .B2(b[21]), .A(n1877), .ZN(n1878) );
  NAND3_X1 U2289 ( .A1(n1880), .A2(n1879), .A3(n1878), .ZN(n1891) );
  NAND2_X1 U2290 ( .A1(n1891), .A2(n1992), .ZN(n1888) );
  NAND2_X1 U2291 ( .A1(n1881), .A2(n2165), .ZN(n1882) );
  OAI21_X1 U2292 ( .B1(n1883), .B2(n2165), .A(n1882), .ZN(n1885) );
  NOR2_X1 U2293 ( .A1(n1885), .A2(n1884), .ZN(n1890) );
  INV_X1 U2294 ( .A(n1891), .ZN(n1887) );
  AOI22_X1 U2295 ( .A1(n1888), .A2(n1890), .B1(n1887), .B2(n1886), .ZN(n2010)
         );
  XNOR2_X1 U2296 ( .A(n1889), .B(n2010), .ZN(\intadd_58/A[3] ) );
  XNOR2_X1 U2297 ( .A(n1890), .B(n1992), .ZN(n1892) );
  XNOR2_X1 U2298 ( .A(n1892), .B(n1891), .ZN(\intadd_58/A[2] ) );
  AND2_X1 U2299 ( .A1(n1893), .A2(b[21]), .ZN(n1898) );
  NOR2_X1 U2300 ( .A1(n1994), .A2(b[21]), .ZN(n1897) );
  NAND2_X1 U2301 ( .A1(n1999), .A2(b[20]), .ZN(n1894) );
  OAI21_X1 U2302 ( .B1(n1895), .B2(b[20]), .A(n1894), .ZN(n1896) );
  NOR3_X1 U2303 ( .A1(n1898), .A2(n1897), .A3(n1896), .ZN(\intadd_58/B[1] ) );
  AND2_X1 U2304 ( .A1(a[23]), .A2(b[18]), .ZN(\intadd_58/B[0] ) );
  NOR2_X1 U2305 ( .A1(n1899), .A2(b[23]), .ZN(n1901) );
  AOI211_X1 U2306 ( .C1(b[23]), .C2(n1902), .A(n1901), .B(n1900), .ZN(
        \intadd_58/CI ) );
  XOR2_X1 U2307 ( .A(\intadd_76/SUM[2] ), .B(n1903), .Z(n1908) );
  OAI21_X1 U2309 ( .B1(n1907), .B2(n1906), .A(n1905), .ZN(n1980) );
  MUX2_X1 U2310 ( .A(n1909), .B(n1908), .S(n1980), .Z(\d[18] ) );
  NOR3_X1 U2311 ( .A1(n1912), .A2(n1978), .A3(n1911), .ZN(n1914) );
  NOR2_X1 U2312 ( .A1(n1914), .A2(n1913), .ZN(\intadd_57/CI ) );
  NOR2_X1 U2313 ( .A1(n1947), .A2(n1915), .ZN(n1950) );
  NAND3_X1 U2314 ( .A1(n1917), .A2(n1933), .A3(n1916), .ZN(n1918) );
  NOR2_X1 U2315 ( .A1(n1919), .A2(n1918), .ZN(n1928) );
  NAND2_X1 U2316 ( .A1(n1922), .A2(n1921), .ZN(n1923) );
  NAND3_X1 U2317 ( .A1(n1925), .A2(n1924), .A3(n1923), .ZN(n1926) );
  AOI22_X1 U2318 ( .A1(n1929), .A2(n1928), .B1(n1927), .B2(n1926), .ZN(n2148)
         );
  NOR2_X1 U2319 ( .A1(n1930), .A2(n1937), .ZN(n1931) );
  XOR2_X1 U2320 ( .A(n2148), .B(n1931), .Z(\d[38]_BAR ) );
  XOR2_X1 U2321 ( .A(\intadd_53/SUM[4] ), .B(n1949), .Z(n1932) );
  XNOR2_X1 U2322 ( .A(n1950), .B(n1932), .ZN(\d[25] ) );
  AOI21_X1 U2323 ( .B1(n1986), .B2(n1933), .A(n1987), .ZN(n2126) );
  NOR2_X1 U2324 ( .A1(n2125), .A2(n2122), .ZN(n1934) );
  XOR2_X1 U2325 ( .A(n2126), .B(n1934), .Z(\d[36]_BAR ) );
  XOR2_X1 U2326 ( .A(n1936), .B(n1935), .Z(\d[2] ) );
  OAI21_X1 U2327 ( .B1(n1938), .B2(n1937), .A(n2024), .ZN(n1941) );
  INV_X1 U2328 ( .A(n2025), .ZN(n1939) );
  NAND2_X1 U2329 ( .A1(n1939), .A2(n2130), .ZN(n1940) );
  XNOR2_X1 U2330 ( .A(n1941), .B(n1940), .ZN(\d[39]_BAR ) );
  INV_X1 U2331 ( .A(n1942), .ZN(n1943) );
  NOR3_X1 U2332 ( .A1(\intadd_56/n1 ), .A2(n1944), .A3(n1943), .ZN(n1945) );
  NOR3_X1 U2333 ( .A1(n1947), .A2(n1946), .A3(n1945), .ZN(n1948) );
  OAI22_X1 U2334 ( .A1(n1950), .A2(n1949), .B1(n1948), .B2(\intadd_53/SUM[4] ), 
        .ZN(n2065) );
  AOI21_X1 U2335 ( .B1(n2065), .B2(n1952), .A(n1951), .ZN(n2100) );
  NAND2_X1 U2336 ( .A1(n2100), .A2(n1953), .ZN(n1964) );
  INV_X1 U2337 ( .A(n2107), .ZN(n1958) );
  AOI21_X1 U2338 ( .B1(\intadd_51/B[4] ), .B2(\intadd_51/A[4] ), .A(n1954), 
        .ZN(n1955) );
  OAI21_X1 U2339 ( .B1(n1966), .B2(n1955), .A(n2018), .ZN(n2074) );
  AOI211_X1 U2340 ( .C1(n2101), .C2(n2107), .A(n1956), .B(n2074), .ZN(n1957)
         );
  OAI21_X1 U2341 ( .B1(n1964), .B2(n1958), .A(n1957), .ZN(n1959) );
  NAND2_X1 U2342 ( .A1(n1959), .A2(n2104), .ZN(n1962) );
  NAND2_X1 U2343 ( .A1(n2076), .A2(n2078), .ZN(n1961) );
  XNOR2_X1 U2344 ( .A(n1962), .B(n1961), .ZN(\d[32] ) );
  NAND2_X1 U2345 ( .A1(n1964), .A2(n1963), .ZN(n2075) );
  NAND2_X1 U2346 ( .A1(n2017), .A2(n1966), .ZN(n1967) );
  XOR2_X1 U2347 ( .A(n2075), .B(n1967), .Z(\d[29] ) );
  NOR2_X1 U2348 ( .A1(n2043), .A2(n1968), .ZN(n2048) );
  NOR2_X1 U2349 ( .A1(n2045), .A2(n2047), .ZN(n1969) );
  XOR2_X1 U2350 ( .A(n2048), .B(n1969), .Z(\d[3] ) );
  NAND2_X1 U2351 ( .A1(n1971), .A2(n1970), .ZN(n1973) );
  XNOR2_X1 U2352 ( .A(n1973), .B(n1972), .ZN(n1974) );
  XOR2_X1 U2353 ( .A(\intadd_72/SUM[0] ), .B(n1974), .Z(\d[5]_BAR ) );
  AND2_X1 U2354 ( .A1(n1975), .A2(n2051), .ZN(n1976) );
  OAI22_X1 U2355 ( .A1(n2052), .A2(n1977), .B1(\intadd_72/n1 ), .B2(n1976), 
        .ZN(\d[8]_BAR ) );
  AOI21_X1 U2356 ( .B1(n1980), .B2(n1979), .A(n1978), .ZN(n1984) );
  NAND2_X1 U2357 ( .A1(n1982), .A2(n1981), .ZN(n1983) );
  XNOR2_X1 U2358 ( .A(n1984), .B(n1983), .ZN(\d[19] ) );
  NAND2_X1 U2360 ( .A1(n1986), .A2(n1985), .ZN(n1990) );
  NOR2_X1 U2361 ( .A1(n1988), .A2(n1987), .ZN(n1989) );
  XNOR2_X1 U2362 ( .A(n1990), .B(n1989), .ZN(\d[35] ) );
  NOR2_X1 U2363 ( .A1(n1992), .A2(n1991), .ZN(n2000) );
  NOR2_X1 U2364 ( .A1(n2167), .A2(a[22]), .ZN(n1997) );
  NAND2_X1 U2365 ( .A1(n1997), .A2(n2165), .ZN(n1993) );
  NAND2_X1 U2366 ( .A1(n1994), .A2(n1993), .ZN(n2005) );
  OAI211_X1 U2367 ( .C1(n1995), .C2(n2000), .A(n2005), .B(n1998), .ZN(n2164)
         );
  NAND3_X1 U2368 ( .A1(n1998), .A2(n1997), .A3(n1996), .ZN(n2003) );
  NAND2_X1 U2369 ( .A1(n1999), .A2(b[23]), .ZN(n2002) );
  NAND3_X1 U2370 ( .A1(n2003), .A2(n2002), .A3(n2001), .ZN(n2004) );
  NOR2_X1 U2371 ( .A1(n2005), .A2(n2004), .ZN(n2161) );
  NAND2_X1 U2373 ( .A1(a[23]), .A2(b[22]), .ZN(n2163) );
  NAND2_X1 U2375 ( .A1(n2010), .A2(n2009), .ZN(n2014) );
  INV_X1 U2376 ( .A(n2010), .ZN(n2011) );
  AOI22_X1 U2377 ( .A1(n2014), .A2(n2013), .B1(n2012), .B2(n2011), .ZN(n2175)
         );
  XOR2_X1 U2378 ( .A(n2171), .B(n2175), .Z(n2015) );
  XNOR2_X1 U2379 ( .A(\intadd_58/n1 ), .B(n2015), .ZN(\d[46]_BAR ) );
  NAND2_X1 U2380 ( .A1(n1964), .A2(n2016), .ZN(n2108) );
  NAND2_X1 U2381 ( .A1(n2108), .A2(n2017), .ZN(n2022) );
  INV_X1 U2382 ( .A(n2018), .ZN(n2020) );
  NOR2_X1 U2383 ( .A1(n2020), .A2(n2019), .ZN(n2021) );
  XOR2_X1 U2384 ( .A(n2022), .B(n2021), .Z(\d[30] ) );
  NAND2_X1 U2385 ( .A1(n2148), .A2(n2023), .ZN(n2132) );
  NOR2_X1 U2386 ( .A1(n2025), .A2(n2024), .ZN(n2129) );
  NOR2_X1 U2387 ( .A1(n2026), .A2(n2129), .ZN(n2145) );
  NAND2_X1 U2388 ( .A1(n2132), .A2(n2145), .ZN(n2139) );
  INV_X1 U2389 ( .A(n2032), .ZN(n2134) );
  INV_X1 U2390 ( .A(n2027), .ZN(n2028) );
  NAND2_X1 U2391 ( .A1(n2028), .A2(n2036), .ZN(n2030) );
  AOI21_X1 U2392 ( .B1(n2139), .B2(n2134), .A(n2030), .ZN(n2035) );
  NOR2_X1 U2393 ( .A1(n2148), .A2(n2029), .ZN(n2038) );
  INV_X1 U2394 ( .A(n2030), .ZN(n2031) );
  NOR4_X1 U2395 ( .A1(n2038), .A2(n2033), .A3(n2032), .A4(n2031), .ZN(n2034)
         );
  OAI21_X1 U2396 ( .B1(n2038), .B2(n2037), .A(n2036), .ZN(n2042) );
  INV_X1 U2397 ( .A(n2140), .ZN(n2040) );
  NAND2_X1 U2398 ( .A1(n2040), .A2(n2039), .ZN(n2041) );
  XNOR2_X1 U2399 ( .A(n2042), .B(n2041), .ZN(\d[42]_BAR ) );
  XOR2_X1 U2400 ( .A(n2044), .B(n2043), .Z(n2050) );
  INV_X1 U2401 ( .A(n2045), .ZN(n2046) );
  OAI21_X1 U2402 ( .B1(n2048), .B2(n2047), .A(n2046), .ZN(n2049) );
  XOR2_X1 U2403 ( .A(n2050), .B(n2049), .Z(\d[4]_BAR ) );
  NAND2_X1 U2404 ( .A1(n2052), .A2(n2051), .ZN(n2056) );
  NAND2_X1 U2405 ( .A1(n2054), .A2(n2053), .ZN(n2055) );
  XOR2_X1 U2406 ( .A(n2056), .B(n2055), .Z(\d[9]_BAR ) );
  XNOR2_X1 U2407 ( .A(n2092), .B(\intadd_64/n1 ), .ZN(n2061) );
  INV_X1 U2408 ( .A(n2057), .ZN(n2090) );
  INV_X1 U2409 ( .A(n2060), .ZN(n2089) );
  NOR3_X1 U2410 ( .A1(n2092), .A2(n2089), .A3(\intadd_64/n1 ), .ZN(n2058) );
  AOI21_X1 U2411 ( .B1(n2092), .B2(n2090), .A(n2058), .ZN(n2059) );
  OAI21_X1 U2412 ( .B1(n2061), .B2(n2060), .A(n2059), .ZN(\d[15]_BAR ) );
  XOR2_X1 U2413 ( .A(n2063), .B(n2062), .Z(n2064) );
  XNOR2_X1 U2414 ( .A(\intadd_57/n1 ), .B(n2064), .ZN(\d[24]_BAR ) );
  XOR2_X1 U2415 ( .A(\intadd_52/SUM[4] ), .B(\intadd_53/n1 ), .Z(n2066) );
  INV_X1 U2416 ( .A(n2066), .ZN(n2067) );
  MUX2_X1 U2417 ( .A(n2067), .B(n2066), .S(n2065), .Z(\d[26]_BAR ) );
  OAI21_X1 U2418 ( .B1(n2065), .B2(n2069), .A(n2068), .ZN(n2073) );
  NAND2_X1 U2419 ( .A1(n2071), .A2(n2070), .ZN(n2072) );
  XNOR2_X1 U2420 ( .A(n2073), .B(n2072), .ZN(\d[27]_BAR ) );
  AOI21_X1 U2421 ( .B1(n2075), .B2(n2107), .A(n2074), .ZN(n2102) );
  OAI21_X1 U2422 ( .B1(n2102), .B2(n2106), .A(n2077), .ZN(n2113) );
  NAND2_X1 U2423 ( .A1(n2113), .A2(n2078), .ZN(n2081) );
  NOR2_X1 U2424 ( .A1(n2111), .A2(n2079), .ZN(n2080) );
  XNOR2_X1 U2425 ( .A(n2081), .B(n2080), .ZN(\d[33]_BAR ) );
  AOI21_X1 U2427 ( .B1(a[0]), .B2(n2084), .A(n2083), .ZN(n2087) );
  OAI22_X1 U2428 ( .A1(n2087), .A2(n2086), .B1(n2085), .B2(n2084), .ZN(\d[1] )
         );
  AOI21_X1 U2430 ( .B1(n2092), .B2(n2091), .A(n2090), .ZN(n2097) );
  INV_X1 U2431 ( .A(n2093), .ZN(n2095) );
  NAND2_X1 U2432 ( .A1(n2095), .A2(n2094), .ZN(n2096) );
  XNOR2_X1 U2433 ( .A(n2097), .B(n2096), .ZN(\d[16] ) );
  NOR2_X1 U2434 ( .A1(n2101), .A2(n2098), .ZN(n2099) );
  OAI22_X1 U2435 ( .A1(n1964), .A2(n2101), .B1(n2100), .B2(n2099), .ZN(\d[28] ) );
  AOI21_X1 U2436 ( .B1(n2104), .B2(n2103), .A(n2102), .ZN(n2110) );
  AOI211_X1 U2437 ( .C1(n2108), .C2(n2107), .A(n2106), .B(n2105), .ZN(n2109)
         );
  NOR2_X1 U2438 ( .A1(n2110), .A2(n2109), .ZN(\d[31] ) );
  AOI21_X1 U2439 ( .B1(n2113), .B2(n2112), .A(n2111), .ZN(n2117) );
  NOR2_X1 U2440 ( .A1(n2115), .A2(n2114), .ZN(n2116) );
  XOR2_X1 U2441 ( .A(n2117), .B(n2116), .Z(\d[34] ) );
  XNOR2_X1 U2442 ( .A(\intadd_59/n1 ), .B(n2118), .ZN(n2121) );
  OAI211_X1 U2444 ( .C1(n2120), .C2(n2122), .A(n2121), .B(n2119), .ZN(n2128)
         );
  INV_X1 U2445 ( .A(n2121), .ZN(n2124) );
  OAI211_X1 U2446 ( .C1(n2126), .C2(n2125), .A(n2124), .B(n2123), .ZN(n2127)
         );
  NAND2_X1 U2447 ( .A1(n2128), .A2(n2127), .ZN(\d[37]_BAR ) );
  INV_X1 U2448 ( .A(n2129), .ZN(n2131) );
  NAND3_X1 U2449 ( .A1(n2132), .A2(n2131), .A3(n2130), .ZN(n2136) );
  NAND2_X1 U2450 ( .A1(n2134), .A2(n2133), .ZN(n2135) );
  XOR2_X1 U2451 ( .A(n2136), .B(n2135), .Z(\d[40] ) );
  AOI21_X1 U2452 ( .B1(n2139), .B2(n2138), .A(n2137), .ZN(n2141) );
  NOR2_X1 U2453 ( .A1(n2141), .A2(n2140), .ZN(n2144) );
  NOR2_X1 U2454 ( .A1(n2152), .A2(n2142), .ZN(n2143) );
  XNOR2_X1 U2455 ( .A(n2144), .B(n2143), .ZN(\d[43] ) );
  OAI21_X1 U2456 ( .B1(n2148), .B2(n2147), .A(n2146), .ZN(n2151) );
  AOI21_X1 U2457 ( .B1(n2151), .B2(n2150), .A(n2149), .ZN(n2155) );
  NOR2_X1 U2458 ( .A1(n2155), .A2(n2152), .ZN(n2156) );
  AOI21_X1 U2459 ( .B1(n2157), .B2(n2153), .A(n2156), .ZN(n2160) );
  NOR2_X1 U2460 ( .A1(n2155), .A2(n2154), .ZN(n2159) );
  OAI22_X1 U2461 ( .A1(n2160), .A2(n2159), .B1(n2158), .B2(n2157), .ZN(\d[44] ) );
  INV_X1 U2462 ( .A(n2171), .ZN(n2173) );
  NAND2_X1 U2463 ( .A1(n2161), .A2(n2163), .ZN(n2162) );
  OAI21_X1 U2464 ( .B1(n2164), .B2(n2163), .A(n2162), .ZN(n2170) );
  XOR2_X1 U2465 ( .A(n2166), .B(n2165), .Z(n2168) );
  NOR2_X1 U2466 ( .A1(n2168), .A2(n2167), .ZN(n2169) );
  XNOR2_X1 U2467 ( .A(n2170), .B(n2169), .ZN(n2172) );
  INV_X1 U2468 ( .A(n2172), .ZN(n2174) );
  AOI21_X1 U2469 ( .B1(n2175), .B2(n2173), .A(n2174), .ZN(n2181) );
  OAI21_X1 U2470 ( .B1(n2175), .B2(n2173), .A(n2174), .ZN(n2179) );
  NAND2_X1 U2471 ( .A1(n2172), .A2(n2171), .ZN(n2177) );
  NAND2_X1 U2472 ( .A1(n2174), .A2(n2173), .ZN(n2176) );
  MUX2_X1 U2473 ( .A(n2177), .B(n2176), .S(n2175), .Z(n2178) );
  OAI21_X1 U2474 ( .B1(\intadd_58/n1 ), .B2(n2179), .A(n2178), .ZN(n2180) );
  AOI21_X1 U2475 ( .B1(\intadd_58/n1 ), .B2(n2181), .A(n2180), .ZN(\d[47] ) );
  INV_X1 U1 ( .A(b[0]), .ZN(n2084) );
  AND2_X1 U2 ( .A1(a[0]), .A2(b[0]), .ZN(\d[0] ) );
  INV_X1 U3 ( .A(n2119), .ZN(n2125) );
  NAND2_X1 U6 ( .A1(\intadd_59/SUM[3] ), .A2(\intadd_48/n1 ), .ZN(n2119) );
  OR2_X2 U7 ( .A1(n2060), .A2(\intadd_64/n1 ), .ZN(n2091) );
  INV_X1 U11 ( .A(n1985), .ZN(n2115) );
  NAND2_X1 U12 ( .A1(\intadd_47/SUM[4] ), .A2(\intadd_49/n1 ), .ZN(n1985) );
  INV_X1 U15 ( .A(n1906), .ZN(n1904) );
  NOR2_X1 U17 ( .A1(\intadd_66/n1 ), .A2(\intadd_65/SUM[3] ), .ZN(n1906) );
  INV_X1 U18 ( .A(n2101), .ZN(n1963) );
  NOR2_X1 U22 ( .A1(n572), .A2(n573), .ZN(n2101) );
  XOR2_X1 U23 ( .A(n2163), .B(n2199), .Z(n2171) );
  NAND2_X1 U24 ( .A1(n2006), .A2(n2164), .ZN(n2199) );
  INV_X1 U28 ( .A(n1978), .ZN(n1910) );
  NOR2_X1 U35 ( .A1(n1903), .A2(\intadd_76/SUM[2] ), .ZN(n1978) );
  NAND3_X1 U37 ( .A1(n1925), .A2(n594), .A3(n2200), .ZN(n1986) );
  NAND3_X1 U42 ( .A1(n1947), .A2(n1917), .A3(n593), .ZN(n2200) );
  INV_X1 U43 ( .A(n578), .ZN(n2016) );
  NAND2_X1 U46 ( .A1(n1963), .A2(n1966), .ZN(n578) );
  NOR3_X1 U50 ( .A1(n2201), .A2(n2111), .A3(n2105), .ZN(n586) );
  INV_X1 U51 ( .A(n2076), .ZN(n2201) );
  NAND2_X1 U60 ( .A1(n381), .A2(n1920), .ZN(n2076) );
  INV_X1 U61 ( .A(n327), .ZN(n326) );
  OAI22_X1 U63 ( .A1(n308), .A2(n309), .B1(n307), .B2(n2203), .ZN(n327) );
  INV_X1 U66 ( .A(n312), .ZN(n2203) );
  INV_X1 U69 ( .A(n1913), .ZN(n1982) );
  NOR2_X1 U72 ( .A1(n353), .A2(\intadd_77/SUM[2] ), .ZN(n1913) );
  AOI21_X1 U73 ( .B1(n580), .B2(n582), .A(n2204), .ZN(n1920) );
  INV_X1 U74 ( .A(\intadd_50/SUM[4] ), .ZN(n2204) );
  AOI22_X1 U75 ( .A1(\intadd_53/SUM[3] ), .A2(\intadd_52/SUM[2] ), .B1(n569), 
        .B2(n2205), .ZN(n1946) );
  OR2_X1 U78 ( .A1(\intadd_53/SUM[3] ), .A2(\intadd_52/SUM[2] ), .ZN(n2205) );
  OAI211_X1 U80 ( .C1(b[19]), .C2(b[18]), .A(a[23]), .B(n2206), .ZN(n319) );
  NAND2_X1 U82 ( .A1(b[19]), .A2(b[18]), .ZN(n2206) );
  OAI21_X1 U84 ( .B1(\intadd_62/n1 ), .B2(n563), .A(n2207), .ZN(n572) );
  INV_X1 U86 ( .A(n2208), .ZN(n2207) );
  AOI21_X1 U87 ( .B1(\intadd_62/n1 ), .B2(n563), .A(n564), .ZN(n2208) );
  OAI21_X1 U89 ( .B1(n357), .B2(n356), .A(n2209), .ZN(\intadd_57/A[1] ) );
  INV_X1 U90 ( .A(n2209), .ZN(n114) );
  NAND2_X1 U92 ( .A1(\intadd_67/n1 ), .A2(\intadd_55/SUM[3] ), .ZN(n2209) );
  AOI21_X1 U93 ( .B1(\intadd_79/n1 ), .B2(\intadd_52/SUM[1] ), .A(n2210), .ZN(
        n179) );
  OAI21_X1 U94 ( .B1(\intadd_79/n1 ), .B2(\intadd_52/SUM[1] ), .A(n368), .ZN(
        n2210) );
  OR3_X1 U95 ( .A1(\intadd_66/SUM[3] ), .A2(n340), .A3(\intadd_64/n1 ), .ZN(
        n338) );
  OAI211_X1 U96 ( .C1(b[17]), .C2(b[16]), .A(a[23]), .B(n2211), .ZN(n300) );
  NAND2_X1 U97 ( .A1(b[17]), .A2(b[16]), .ZN(n2211) );
  OAI211_X1 U99 ( .C1(b[13]), .C2(b[12]), .A(a[23]), .B(n2212), .ZN(n866) );
  NAND2_X1 U101 ( .A1(b[13]), .A2(b[12]), .ZN(n2212) );
  INV_X1 U102 ( .A(b[17]), .ZN(n893) );
  INV_X1 U103 ( .A(b[16]), .ZN(n1246) );
  NAND2_X1 U105 ( .A1(b[17]), .A2(b[16]), .ZN(n268) );
  INV_X1 U106 ( .A(\intadd_65/SUM[1] ), .ZN(n341) );
  OAI21_X1 U107 ( .B1(\intadd_66/SUM[2] ), .B2(\intadd_75/n1 ), .A(n2213), 
        .ZN(n343) );
  AOI21_X1 U109 ( .B1(\intadd_66/SUM[2] ), .B2(\intadd_75/n1 ), .A(
        \intadd_65/SUM[1] ), .ZN(n2213) );
  INV_X1 U110 ( .A(n581), .ZN(n381) );
  NOR2_X1 U114 ( .A1(\intadd_71/SUM[2] ), .A2(\intadd_50/SUM[3] ), .ZN(n581)
         );
  AOI21_X1 U116 ( .B1(b[11]), .B2(b[10]), .A(n2214), .ZN(n253) );
  INV_X1 U118 ( .A(n916), .ZN(n2214) );
  NOR2_X1 U123 ( .A1(n219), .A2(n218), .ZN(n916) );
  OAI211_X1 U124 ( .C1(b[9]), .C2(b[8]), .A(a[23]), .B(n2215), .ZN(n993) );
  NAND2_X1 U125 ( .A1(b[9]), .A2(b[8]), .ZN(n2215) );
  INV_X1 U136 ( .A(n1525), .ZN(n1524) );
  NAND2_X1 U140 ( .A1(n1527), .A2(n1526), .ZN(n1525) );
  INV_X1 U144 ( .A(n1145), .ZN(n1152) );
  NAND2_X1 U152 ( .A1(n1143), .A2(n1144), .ZN(n1145) );
  INV_X1 U153 ( .A(n1461), .ZN(n1501) );
  NAND2_X1 U154 ( .A1(n1455), .A2(n1456), .ZN(n1461) );
  OR2_X2 U156 ( .A1(n1628), .A2(n1627), .ZN(n1658) );
  XOR2_X1 U162 ( .A(n523), .B(n525), .Z(n526) );
  XNOR2_X1 U163 ( .A(n435), .B(n457), .ZN(n525) );
  AOI21_X1 U164 ( .B1(n1711), .B2(b[10]), .A(n2216), .ZN(n1632) );
  OAI22_X1 U168 ( .A1(b[10]), .A2(n2217), .B1(n1510), .B2(n1511), .ZN(n2216)
         );
  INV_X1 U170 ( .A(n1712), .ZN(n2217) );
  OAI21_X1 U173 ( .B1(b[21]), .B2(n1856), .A(n2218), .ZN(n1464) );
  AOI22_X1 U175 ( .A1(n1309), .A2(n1867), .B1(b[21]), .B2(n2219), .ZN(n2218)
         );
  INV_X1 U176 ( .A(n1855), .ZN(n2219) );
  OAI21_X1 U177 ( .B1(b[10]), .B2(n1697), .A(n2220), .ZN(n1592) );
  AOI22_X1 U179 ( .A1(n1505), .A2(n1506), .B1(b[10]), .B2(n2221), .ZN(n2220)
         );
  INV_X1 U183 ( .A(n1698), .ZN(n2221) );
  INV_X1 U184 ( .A(n1380), .ZN(n1379) );
  AOI211_X1 U196 ( .C1(b[1]), .C2(n190), .A(n2009), .B(b[0]), .ZN(n1380) );
  NOR3_X1 U201 ( .A1(n232), .A2(b[23]), .A3(a[12]), .ZN(n183) );
  AOI211_X1 U208 ( .C1(n1742), .C2(b[10]), .A(n1399), .B(n2222), .ZN(n1576) );
  INV_X1 U211 ( .A(n2223), .ZN(n2222) );
  MUX2_X1 U224 ( .A(n1698), .B(n1697), .S(b[11]), .Z(n2223) );
  INV_X1 U229 ( .A(n1413), .ZN(n1395) );
  NAND2_X1 U230 ( .A1(n735), .A2(n736), .ZN(n1413) );
  INV_X1 U231 ( .A(n2224), .ZN(n1527) );
  OAI21_X1 U237 ( .B1(n2084), .B2(n1453), .A(\intadd_58/A[1] ), .ZN(n2224) );
  NOR2_X1 U247 ( .A1(n1443), .A2(n1442), .ZN(\intadd_58/A[1] ) );
  AND2_X2 U249 ( .A1(n1478), .A2(b[3]), .ZN(n1582) );
  OAI21_X1 U251 ( .B1(b[23]), .B2(n1856), .A(n2225), .ZN(n1368) );
  AOI22_X1 U254 ( .A1(n1996), .A2(n1867), .B1(b[23]), .B2(n2226), .ZN(n2225)
         );
  INV_X1 U260 ( .A(n1855), .ZN(n2226) );
  OAI21_X1 U268 ( .B1(b[17]), .B2(n1856), .A(n2227), .ZN(n1566) );
  AOI22_X1 U272 ( .A1(n1246), .A2(n1867), .B1(b[17]), .B2(n2228), .ZN(n2227)
         );
  INV_X1 U275 ( .A(n1855), .ZN(n2228) );
  INV_X1 U283 ( .A(n1647), .ZN(n628) );
  NAND2_X1 U284 ( .A1(n621), .A2(n622), .ZN(n1647) );
  OAI21_X1 U286 ( .B1(b[15]), .B2(n1856), .A(n2230), .ZN(n1662) );
  AOI22_X1 U295 ( .A1(n1602), .A2(n1867), .B1(b[15]), .B2(n2231), .ZN(n2230)
         );
  INV_X1 U299 ( .A(n1855), .ZN(n2231) );
  OAI21_X1 U307 ( .B1(b[18]), .B2(n1856), .A(n2232), .ZN(n1534) );
  AOI22_X1 U310 ( .A1(n893), .A2(n1867), .B1(b[18]), .B2(n2233), .ZN(n2232) );
  INV_X1 U312 ( .A(n1855), .ZN(n2233) );
  OR2_X2 U315 ( .A1(n457), .A2(n456), .ZN(n459) );
  OR2_X2 U320 ( .A1(n519), .A2(n518), .ZN(n521) );
  NOR3_X1 U323 ( .A1(n1250), .A2(b[23]), .A3(a[8]), .ZN(n970) );
  INV_X1 U333 ( .A(n101), .ZN(n2234) );
  INV_X1 U334 ( .A(n1843), .ZN(n2235) );
  OAI22_X2 U335 ( .A1(n2235), .A2(n2234), .B1(n1842), .B2(\intadd_46/SUM[0] ), 
        .ZN(n109) );
  INV_X1 U343 ( .A(n770), .ZN(n293) );
  NAND2_X1 U346 ( .A1(a[17]), .A2(n783), .ZN(n770) );
  INV_X1 U349 ( .A(n1623), .ZN(n1652) );
  AOI211_X1 U350 ( .C1(n1611), .C2(n1689), .A(n1613), .B(n1612), .ZN(n1623) );
  INV_X1 U351 ( .A(n762), .ZN(n759) );
  NAND2_X1 U362 ( .A1(n753), .A2(n754), .ZN(n762) );
  INV_X1 U364 ( .A(n1187), .ZN(n1135) );
  NOR2_X1 U365 ( .A1(n1999), .A2(n1869), .ZN(n1187) );
  AOI21_X1 U366 ( .B1(a[23]), .B2(b[7]), .A(n2236), .ZN(n615) );
  INV_X1 U381 ( .A(n1030), .ZN(n2236) );
  NAND2_X1 U382 ( .A1(b[6]), .A2(a[23]), .ZN(n1030) );
  OAI21_X1 U383 ( .B1(b[19]), .B2(n1856), .A(n2238), .ZN(n735) );
  AOI22_X1 U408 ( .A1(n1247), .A2(n1867), .B1(b[19]), .B2(n2239), .ZN(n2238)
         );
  INV_X1 U430 ( .A(n1855), .ZN(n2239) );
  INV_X1 U433 ( .A(n159), .ZN(n158) );
  NAND2_X1 U434 ( .A1(a[19]), .A2(a[20]), .ZN(n159) );
  INV_X1 U448 ( .A(n1895), .ZN(n1869) );
  NAND2_X1 U449 ( .A1(a[23]), .A2(n438), .ZN(n1895) );
  INV_X1 U454 ( .A(n61), .ZN(n1835) );
  NAND2_X1 U455 ( .A1(n53), .A2(n54), .ZN(n61) );
  AND2_X1 U456 ( .A1(n70), .A2(n2240), .ZN(n80) );
  XNOR2_X1 U460 ( .A(n74), .B(n73), .ZN(n2240) );
  INV_X1 U461 ( .A(n1448), .ZN(n989) );
  NAND2_X1 U462 ( .A1(n1442), .A2(n1517), .ZN(n1448) );
  NOR2_X1 U471 ( .A1(a[15]), .A2(n627), .ZN(n1478) );
  INV_X1 U477 ( .A(n1730), .ZN(n883) );
  NAND2_X1 U482 ( .A1(a[11]), .A2(n123), .ZN(n1730) );
  AOI211_X1 U516 ( .C1(b[0]), .C2(n2242), .A(\intadd_54/A[0] ), .B(n2241), 
        .ZN(n1816) );
  NOR2_X1 U517 ( .A1(b[0]), .A2(n1775), .ZN(n2241) );
  INV_X1 U540 ( .A(n1774), .ZN(n2242) );
  INV_X1 U541 ( .A(n1530), .ZN(n1434) );
  NOR2_X1 U555 ( .A1(a[17]), .A2(n783), .ZN(n1530) );
  INV_X1 U556 ( .A(n1726), .ZN(n1702) );
  NOR2_X1 U558 ( .A1(n124), .A2(n125), .ZN(n1726) );
  NOR3_X1 U559 ( .A1(n2243), .A2(n649), .A3(a[13]), .ZN(n1389) );
  INV_X1 U564 ( .A(n1706), .ZN(n2243) );
  NAND2_X1 U565 ( .A1(a[12]), .A2(a[11]), .ZN(n1706) );
  NOR3_X1 U566 ( .A1(n2244), .A2(a[17]), .A3(n213), .ZN(n1529) );
  INV_X1 U579 ( .A(n783), .ZN(n2244) );
  NAND2_X1 U580 ( .A1(a[16]), .A2(a[15]), .ZN(n783) );
  INV_X1 U590 ( .A(n1836), .ZN(n60) );
  NAND2_X1 U591 ( .A1(n55), .A2(n56), .ZN(n1836) );
  INV_X1 U634 ( .A(n2166), .ZN(n1234) );
  NAND2_X1 U638 ( .A1(a[22]), .A2(a[21]), .ZN(n2166) );
  INV_X1 U643 ( .A(n35), .ZN(n1972) );
  OAI22_X1 U644 ( .A1(n27), .A2(n28), .B1(n26), .B2(n2247), .ZN(n35) );
  AOI22_X1 U645 ( .A1(n1805), .A2(n1806), .B1(n87), .B2(n2245), .ZN(n1847) );
  OR2_X1 U660 ( .A1(n1805), .A2(n1806), .ZN(n2245) );
  INV_X1 U707 ( .A(n1810), .ZN(n1809) );
  NAND2_X1 U748 ( .A1(n1783), .A2(n1784), .ZN(n1810) );
  INV_X1 U749 ( .A(n1811), .ZN(n1808) );
  NAND2_X1 U758 ( .A1(n1785), .A2(n1786), .ZN(n1811) );
  INV_X1 U760 ( .A(n31), .ZN(n2247) );
  NAND2_X1 U761 ( .A1(n2084), .A2(n90), .ZN(n70) );
  OAI21_X1 U767 ( .B1(b[9]), .B2(n1856), .A(n2248), .ZN(n1845) );
  AOI22_X1 U768 ( .A1(n1694), .A2(n1867), .B1(b[9]), .B2(n2249), .ZN(n2248) );
  INV_X1 U789 ( .A(n1855), .ZN(n2249) );
  XNOR2_X1 U794 ( .A(a[13]), .B(a[14]), .ZN(n627) );
  INV_X1 U795 ( .A(n117), .ZN(n1443) );
  NAND2_X1 U827 ( .A1(a[18]), .A2(a[17]), .ZN(n117) );
  OAI21_X1 U828 ( .B1(b[6]), .B2(n1856), .A(n2250), .ZN(n1778) );
  AOI22_X1 U871 ( .A1(n1611), .A2(n1867), .B1(b[6]), .B2(n2251), .ZN(n2250) );
  INV_X1 U903 ( .A(n1855), .ZN(n2251) );
  INV_X1 U924 ( .A(n1771), .ZN(n1062) );
  NAND2_X1 U925 ( .A1(a[7]), .A2(n645), .ZN(n1771) );
  OAI21_X1 U1002 ( .B1(b[4]), .B2(n1856), .A(n2252), .ZN(n27) );
  AOI22_X1 U1003 ( .A1(n1787), .A2(n1867), .B1(b[4]), .B2(n2253), .ZN(n2252)
         );
  INV_X1 U1004 ( .A(n1855), .ZN(n2253) );
  AND2_X2 U1007 ( .A1(n22), .A2(n21), .ZN(n2047) );
  INV_X1 U1056 ( .A(n1711), .ZN(n1751) );
  NOR2_X1 U1057 ( .A1(a[7]), .A2(n645), .ZN(n1711) );
  INV_X1 U1058 ( .A(n1698), .ZN(n1739) );
  NAND2_X1 U1060 ( .A1(a[9]), .A2(n1557), .ZN(n1698) );
  OAI21_X1 U1061 ( .B1(b[3]), .B2(n1856), .A(n2254), .ZN(n23) );
  AOI22_X1 U1063 ( .A1(n1740), .A2(n1867), .B1(b[3]), .B2(n2255), .ZN(n2254)
         );
  INV_X1 U1088 ( .A(n1855), .ZN(n2255) );
  INV_X1 U1108 ( .A(n1788), .ZN(n1860) );
  NAND2_X1 U1109 ( .A1(n38), .A2(\intadd_49/B[0] ), .ZN(n1788) );
  INV_X1 U1257 ( .A(n1789), .ZN(n39) );
  NAND2_X1 U1258 ( .A1(a[5]), .A2(n1179), .ZN(n1789) );
  INV_X1 U1259 ( .A(n1851), .ZN(n1765) );
  NAND2_X1 U1260 ( .A1(a[1]), .A2(n1171), .ZN(n1851) );
  INV_X1 U1261 ( .A(n1849), .ZN(n1763) );
  NAND2_X1 U1273 ( .A1(n1331), .A2(n8), .ZN(n1849) );
  INV_X1 U1274 ( .A(n1850), .ZN(n1764) );
  NAND2_X1 U1275 ( .A1(a[3]), .A2(n8), .ZN(n1850) );
  INV_X1 U1313 ( .A(n1855), .ZN(n2083) );
  NAND2_X1 U1315 ( .A1(a[0]), .A2(n1205), .ZN(n1855) );
  INV_X1 U1316 ( .A(n1867), .ZN(n1858) );
  NOR2_X1 U1405 ( .A1(a[0]), .A2(n1205), .ZN(n1867) );
  INV_X1 U1406 ( .A(n1179), .ZN(n38) );
  NOR2_X1 U1516 ( .A1(a[4]), .A2(a[3]), .ZN(n1179) );
endmodule



    module conf_int_mul__noFF__arch_agnos__w_wrapper_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 ( 
        clk, rst, a, b, d__acc, acc__sel, \d[63] , \d[62] , \d[61] , \d[60] , 
        \d[59] , \d[58]_BAR , \d[57] , \d[56] , \d[55] , \d[54] , \d[53] , 
        \d[51] , \d[50] , \d[49] , \d[48] , \d[47] , \d[46] , \d[45] , \d[44] , 
        \d[43] , \d[41] , \d[40] , \d[39] , \d[38] , \d[37] , \d[36] , \d[35] , 
        \d[34] , \d[32] , \d[19] , \d[18] , \d[17] , \d[16] , \d[15] , \d[14] , 
        \d[13] , \d[12] , \d[11] , \d[10] , \d[9] , \d[8] , \d[7] , \d[6] , 
        \d[5] , \d[4] , \d[3] , \d[2] , \d[1] , \d[0] , \d[52]_BAR , 
        \d[42]_BAR , \d[33]_BAR , \d[31]_BAR , \d[30]_BAR , \d[29]_BAR , 
        \d[28]_BAR , \d[27]_BAR , \d[26]_BAR , \d[25]_BAR , \d[24]_BAR , 
        \d[23]_BAR , \d[22]_BAR , \d[21]_BAR , \d[20]_BAR  );
  input [23:0] a;
  input [23:0] b;
  input [63:0] d__acc;
  input clk, rst, acc__sel;
  output \d[63] , \d[62] , \d[61] , \d[60] , \d[59] , \d[58]_BAR , \d[57] ,
         \d[56] , \d[55] , \d[54] , \d[53] , \d[51] , \d[50] , \d[49] ,
         \d[48] , \d[47] , \d[46] , \d[45] , \d[44] , \d[43] , \d[41] ,
         \d[40] , \d[39] , \d[38] , \d[37] , \d[36] , \d[35] , \d[34] ,
         \d[32] , \d[19] , \d[18] , \d[17] , \d[16] , \d[15] , \d[14] ,
         \d[13] , \d[12] , \d[11] , \d[10] , \d[9] , \d[8] , \d[7] , \d[6] ,
         \d[5] , \d[4] , \d[3] , \d[2] , \d[1] , \d[0] , \d[52]_BAR ,
         \d[42]_BAR , \d[33]_BAR , \d[31]_BAR , \d[30]_BAR , \d[29]_BAR ,
         \d[28]_BAR , \d[27]_BAR , \d[26]_BAR , \d[25]_BAR , \d[24]_BAR ,
         \d[23]_BAR , \d[22]_BAR , \d[21]_BAR , \d[20]_BAR ;
  wire   n1, n2, n3, n4, n5, n6, n9, n10, n12, n14, n16, n18, n20, n22, n24,
         n26, n28, n30, n32, n34, n36, n38, n40, n42, n43, n44, n45, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60;
  wire   [63:0] d;
  wire   [47:0] d__apx;
  assign \d[63]  = d[63];
  assign \d[62]  = d[62];
  assign \d[61]  = d[61];
  assign \d[60]  = d[60];
  assign \d[59]  = d[59];
  assign \d[57]  = d[57];
  assign \d[56]  = d[56];
  assign \d[55]  = d[55];
  assign \d[54]  = d[54];
  assign \d[53]  = d[53];
  assign \d[51]  = d[51];
  assign \d[50]  = d[50];
  assign \d[49]  = d[49];
  assign \d[48]  = d[48];
  assign \d[47]  = d[47];
  assign \d[46]  = d[46];
  assign \d[45]  = d[45];
  assign \d[44]  = d[44];
  assign \d[43]  = d[43];
  assign \d[41]  = d[41];
  assign \d[40]  = d[40];
  assign \d[39]  = d[39];
  assign \d[38]  = d[38];
  assign \d[37]  = d[37];
  assign \d[36]  = d[36];
  assign \d[35]  = d[35];
  assign \d[34]  = d[34];
  assign \d[32]  = d[32];
  assign \d[18]  = d[18];
  assign \d[17]  = d[17];
  assign \d[16]  = d[16];
  assign \d[15]  = d[15];
  assign \d[14]  = d[14];
  assign \d[13]  = d[13];
  assign \d[12]  = d[12];
  assign \d[11]  = d[11];
  assign \d[10]  = d[10];
  assign \d[9]  = d[9];
  assign \d[8]  = d[8];
  assign \d[7]  = d[7];
  assign \d[6]  = d[6];
  assign \d[5]  = d[5];
  assign \d[4]  = d[4];
  assign \d[3]  = d[3];
  assign \d[2]  = d[2];
  assign \d[1]  = d[1];
  assign \d[0]  = d[0];

  INV_X1 U1 ( .A(d__apx[7]), .ZN(n2) );
  INV_X1 U2 ( .A(d__apx[10]), .ZN(n3) );
  INV_X1 U3 ( .A(d__apx[12]), .ZN(n4) );
  INV_X1 U4 ( .A(acc__sel), .ZN(n56) );
  LOGIC0_X1 U5 ( .Z(n1) );
  NAND2_X1 U6 ( .A1(d__acc[60]), .A2(acc__sel), .ZN(n6) );
  NAND2_X1 U7 ( .A1(d__apx[44]), .A2(n56), .ZN(n5) );
  NAND2_X1 U8 ( .A1(n6), .A2(n5), .ZN(d[60]) );
  INV_X2 U9 ( .A(d__acc[49]), .ZN(n9) );
  OAI21_X1 U12 ( .B1(n9), .B2(n56), .A(n59), .ZN(d[49]) );
  NOR2_X1 U13 ( .A1(d__apx[6]), .A2(acc__sel), .ZN(n10) );
  AOI21_X1 U14 ( .B1(d__acc[22]), .B2(acc__sel), .A(n10), .ZN(\d[22]_BAR ) );
  NOR2_X1 U15 ( .A1(d__apx[4]), .A2(acc__sel), .ZN(n12) );
  AOI21_X1 U16 ( .B1(d__acc[20]), .B2(acc__sel), .A(n12), .ZN(\d[20]_BAR ) );
  NOR2_X1 U17 ( .A1(d__apx[8]), .A2(acc__sel), .ZN(n14) );
  AOI21_X1 U18 ( .B1(d__acc[24]), .B2(acc__sel), .A(n14), .ZN(\d[24]_BAR ) );
  NOR2_X1 U19 ( .A1(n2), .A2(acc__sel), .ZN(n16) );
  AOI21_X1 U20 ( .B1(d__acc[23]), .B2(acc__sel), .A(n16), .ZN(\d[23]_BAR ) );
  NOR2_X1 U21 ( .A1(d__apx[5]), .A2(acc__sel), .ZN(n18) );
  AOI21_X1 U22 ( .B1(d__acc[21]), .B2(acc__sel), .A(n18), .ZN(\d[21]_BAR ) );
  NOR2_X1 U23 ( .A1(n3), .A2(acc__sel), .ZN(n20) );
  AOI21_X1 U24 ( .B1(d__acc[26]), .B2(acc__sel), .A(n20), .ZN(\d[26]_BAR ) );
  NOR2_X1 U25 ( .A1(d__apx[9]), .A2(acc__sel), .ZN(n22) );
  AOI21_X1 U26 ( .B1(d__acc[25]), .B2(acc__sel), .A(n22), .ZN(\d[25]_BAR ) );
  NOR2_X1 U27 ( .A1(d__apx[11]), .A2(acc__sel), .ZN(n24) );
  AOI21_X1 U28 ( .B1(d__acc[27]), .B2(acc__sel), .A(n24), .ZN(\d[27]_BAR ) );
  NOR2_X1 U29 ( .A1(n4), .A2(acc__sel), .ZN(n26) );
  AOI21_X1 U30 ( .B1(d__acc[28]), .B2(acc__sel), .A(n26), .ZN(\d[28]_BAR ) );
  NOR2_X1 U31 ( .A1(d__apx[14]), .A2(acc__sel), .ZN(n28) );
  AOI21_X1 U32 ( .B1(d__acc[30]), .B2(acc__sel), .A(n28), .ZN(\d[30]_BAR ) );
  NOR2_X1 U33 ( .A1(d__apx[13]), .A2(acc__sel), .ZN(n30) );
  AOI21_X1 U34 ( .B1(d__acc[29]), .B2(acc__sel), .A(n30), .ZN(\d[29]_BAR ) );
  NOR2_X1 U35 ( .A1(d__apx[15]), .A2(acc__sel), .ZN(n32) );
  AOI21_X1 U36 ( .B1(d__acc[31]), .B2(acc__sel), .A(n32), .ZN(\d[31]_BAR ) );
  NOR2_X1 U37 ( .A1(d__apx[17]), .A2(acc__sel), .ZN(n34) );
  AOI21_X1 U38 ( .B1(d__acc[33]), .B2(acc__sel), .A(n34), .ZN(\d[33]_BAR ) );
  NOR2_X1 U39 ( .A1(d__apx[26]), .A2(acc__sel), .ZN(n36) );
  AOI21_X1 U40 ( .B1(d__acc[42]), .B2(acc__sel), .A(n36), .ZN(\d[42]_BAR ) );
  NOR2_X1 U41 ( .A1(d__apx[42]), .A2(acc__sel), .ZN(n38) );
  AOI21_X1 U42 ( .B1(d__acc[58]), .B2(acc__sel), .A(n38), .ZN(\d[58]_BAR ) );
  NOR2_X1 U43 ( .A1(d__apx[36]), .A2(acc__sel), .ZN(n40) );
  AOI21_X1 U44 ( .B1(d__acc[52]), .B2(acc__sel), .A(n40), .ZN(\d[52]_BAR ) );
  MUX2_X1 U45 ( .A(d__apx[16]), .B(d__acc[32]), .S(acc__sel), .Z(d[32]) );
  MUX2_X1 U46 ( .A(d__apx[18]), .B(d__acc[34]), .S(acc__sel), .Z(d[34]) );
  MUX2_X1 U47 ( .A(d__apx[19]), .B(d__acc[35]), .S(acc__sel), .Z(d[35]) );
  MUX2_X1 U48 ( .A(d__apx[20]), .B(d__acc[36]), .S(acc__sel), .Z(d[36]) );
  MUX2_X1 U49 ( .A(d__apx[21]), .B(d__acc[37]), .S(acc__sel), .Z(d[37]) );
  NAND2_X1 U50 ( .A1(d__acc[38]), .A2(acc__sel), .ZN(n42) );
  OAI21_X1 U51 ( .B1(d__apx[22]), .B2(acc__sel), .A(n42), .ZN(d[38]) );
  NAND2_X1 U52 ( .A1(d__acc[39]), .A2(acc__sel), .ZN(n43) );
  OAI21_X1 U53 ( .B1(d__apx[23]), .B2(acc__sel), .A(n43), .ZN(d[39]) );
  NAND2_X1 U54 ( .A1(d__acc[40]), .A2(acc__sel), .ZN(n44) );
  OAI21_X1 U55 ( .B1(d__apx[24]), .B2(acc__sel), .A(n44), .ZN(d[40]) );
  MUX2_X1 U56 ( .A(d__apx[25]), .B(d__acc[41]), .S(acc__sel), .Z(d[41]) );
  NAND2_X1 U57 ( .A1(d__acc[43]), .A2(acc__sel), .ZN(n45) );
  OAI21_X1 U58 ( .B1(acc__sel), .B2(d__apx[27]), .A(n45), .ZN(d[43]) );
  MUX2_X1 U59 ( .A(d__apx[28]), .B(d__acc[44]), .S(acc__sel), .Z(d[44]) );
  MUX2_X1 U60 ( .A(d__apx[29]), .B(d__acc[45]), .S(acc__sel), .Z(d[45]) );
  MUX2_X1 U61 ( .A(d__apx[30]), .B(d__acc[46]), .S(acc__sel), .Z(d[46]) );
  MUX2_X1 U62 ( .A(d__apx[31]), .B(d__acc[47]), .S(acc__sel), .Z(d[47]) );
  MUX2_X1 U63 ( .A(d__apx[32]), .B(d__acc[48]), .S(acc__sel), .Z(d[48]) );
  NAND2_X1 U67 ( .A1(d__acc[51]), .A2(acc__sel), .ZN(n49) );
  NAND2_X1 U68 ( .A1(d__apx[35]), .A2(n56), .ZN(n48) );
  NAND2_X1 U69 ( .A1(n49), .A2(n48), .ZN(d[51]) );
  NAND2_X1 U70 ( .A1(d__acc[53]), .A2(acc__sel), .ZN(n50) );
  OAI21_X1 U71 ( .B1(d__apx[37]), .B2(acc__sel), .A(n50), .ZN(d[53]) );
  NAND2_X1 U72 ( .A1(d__acc[54]), .A2(acc__sel), .ZN(n51) );
  OAI21_X1 U73 ( .B1(d__apx[38]), .B2(acc__sel), .A(n51), .ZN(d[54]) );
  NAND2_X1 U74 ( .A1(d__acc[55]), .A2(acc__sel), .ZN(n52) );
  OAI21_X1 U75 ( .B1(d__apx[39]), .B2(acc__sel), .A(n52), .ZN(d[55]) );
  MUX2_X1 U76 ( .A(d__apx[40]), .B(d__acc[56]), .S(acc__sel), .Z(d[56]) );
  NAND2_X1 U77 ( .A1(d__acc[57]), .A2(acc__sel), .ZN(n53) );
  OAI21_X1 U78 ( .B1(acc__sel), .B2(d__apx[41]), .A(n53), .ZN(d[57]) );
  MUX2_X1 U79 ( .A(d__apx[43]), .B(d__acc[59]), .S(acc__sel), .Z(d[59]) );
  NAND2_X1 U80 ( .A1(d__acc[61]), .A2(acc__sel), .ZN(n54) );
  OAI21_X1 U81 ( .B1(d__apx[45]), .B2(acc__sel), .A(n54), .ZN(d[61]) );
  NAND2_X1 U82 ( .A1(d__acc[62]), .A2(acc__sel), .ZN(n55) );
  OAI21_X1 U83 ( .B1(d__apx[46]), .B2(acc__sel), .A(n55), .ZN(d[62]) );
  NAND2_X1 U84 ( .A1(d__acc[63]), .A2(acc__sel), .ZN(n58) );
  NAND2_X1 U85 ( .A1(d__apx[47]), .A2(n56), .ZN(n57) );
  NAND2_X1 U86 ( .A1(n58), .A2(n57), .ZN(d[63]) );
  AND2_X1 U87 ( .A1(acc__sel), .A2(d__acc[0]), .ZN(d[0]) );
  AND2_X1 U88 ( .A1(acc__sel), .A2(d__acc[1]), .ZN(d[1]) );
  AND2_X1 U89 ( .A1(acc__sel), .A2(d__acc[2]), .ZN(d[2]) );
  AND2_X1 U90 ( .A1(acc__sel), .A2(d__acc[3]), .ZN(d[3]) );
  AND2_X1 U91 ( .A1(acc__sel), .A2(d__acc[4]), .ZN(d[4]) );
  AND2_X1 U92 ( .A1(acc__sel), .A2(d__acc[5]), .ZN(d[5]) );
  AND2_X1 U93 ( .A1(acc__sel), .A2(d__acc[6]), .ZN(d[6]) );
  AND2_X1 U94 ( .A1(acc__sel), .A2(d__acc[7]), .ZN(d[7]) );
  AND2_X1 U95 ( .A1(acc__sel), .A2(d__acc[8]), .ZN(d[8]) );
  AND2_X1 U96 ( .A1(acc__sel), .A2(d__acc[9]), .ZN(d[9]) );
  AND2_X1 U97 ( .A1(acc__sel), .A2(d__acc[10]), .ZN(d[10]) );
  AND2_X1 U98 ( .A1(acc__sel), .A2(d__acc[11]), .ZN(d[11]) );
  AND2_X1 U99 ( .A1(acc__sel), .A2(d__acc[12]), .ZN(d[12]) );
  AND2_X1 U100 ( .A1(acc__sel), .A2(d__acc[13]), .ZN(d[13]) );
  AND2_X1 U101 ( .A1(acc__sel), .A2(d__acc[14]), .ZN(d[14]) );
  AND2_X1 U102 ( .A1(acc__sel), .A2(d__acc[15]), .ZN(d[15]) );
  MUX2_X1 U103 ( .A(d__apx[0]), .B(d__acc[16]), .S(acc__sel), .Z(d[16]) );
  MUX2_X1 U104 ( .A(d__apx[1]), .B(d__acc[17]), .S(acc__sel), .Z(d[17]) );
  MUX2_X1 U105 ( .A(d__apx[2]), .B(d__acc[18]), .S(acc__sel), .Z(d[18]) );
  MUX2_X1 U106 ( .A(d__apx[3]), .B(d__acc[19]), .S(acc__sel), .Z(\d[19] ) );
  OR2_X1 U10 ( .A1(d__apx[33]), .A2(acc__sel), .ZN(n59) );
  conf_int_mul__noFF__arch_agnos_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 mul__inst ( 
        .clk(clk), .rst(n1), .a(a), .b(b), .\d[47] (d__apx[47]), .\d[44] (
        d__apx[44]), .\d[43] (d__apx[43]), .\d[40] (d__apx[40]), .\d[37]_BAR (
        d__apx[37]), .\d[34] (d__apx[34]), .\d[31] (d__apx[31]), .\d[28] (
        d__apx[28]), .\d[16] (d__apx[16]), .\d[1] (d__apx[1]), .\d[0] (
        d__apx[0]), .\d[33]_BAR (d__apx[33]), .\d[27]_BAR (d__apx[27]), 
        .\d[26]_BAR (d__apx[26]), .\d[24]_BAR (d__apx[24]), .\d[23]_BAR (
        d__apx[23]), .\d[15]_BAR (d__apx[15]), .\d[14]_BAR (d__apx[14]), 
        .\d[11]_BAR (d__apx[11]), .\d[9]_BAR (d__apx[9]), .\d[6]_BAR (
        d__apx[6]), .\d[4]_BAR (d__apx[4]), .\d[42]_BAR (d__apx[42]), 
        .\d[41]_BAR (d__apx[41]), .\d[30] (d__apx[30]), .\d[22]_BAR (
        d__apx[22]), .\d[46]_BAR (d__apx[46]), .\d[35] (d__apx[35]), .\d[19] (
        d__apx[19]), .\d[8]_BAR (d__apx[8]), .\d[5]_BAR (d__apx[5]), .\d[3] (
        d__apx[3]), .\d[29] (d__apx[29]), .\d[32] (d__apx[32]), .\d[39]_BAR (
        d__apx[39]), .\d[2] (d__apx[2]), .\d[36]_BAR (d__apx[36]), .\d[25] (
        d__apx[25]), .\d[13]_BAR (d__apx[13]), .\d[38]_BAR (d__apx[38]), 
        .\d[20] (d__apx[20]), .\d[18] (d__apx[18]), .\d[17]_BAR (d__apx[17]), 
        .\d[45]_BAR (d__apx[45]), .\d[21] (d__apx[21]), .\d[12] (d__apx[12]), 
        .\d[10] (d__apx[10]), .\d[7] (d__apx[7]) );
  INV_X1 U11 ( .A(n60), .ZN(d[50]) );
  AOI22_X1 U64 ( .A1(acc__sel), .A2(d__acc[50]), .B1(n56), .B2(d__apx[34]), 
        .ZN(n60) );
endmodule

