library verilog;
use verilog.vl_types.all;
entity INV_X4_func is
    port(
        A               : in     vl_logic;
        ZN              : out    vl_logic
    );
end INV_X4_func;
