


module conf_int_mul__noFF__arch_agnos_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 ( clk, 
        rst, a, b, \d[47] , \d[44] , \d[43] , \d[40] , \d[37]_BAR , \d[34] , 
        \d[31] , \d[28] , \d[16] , \d[1] , \d[0] , \d[33]_BAR , \d[27]_BAR , 
        \d[26]_BAR , \d[24]_BAR , \d[23]_BAR , \d[15]_BAR , \d[14]_BAR , 
        \d[11]_BAR , \d[9]_BAR , \d[4]_BAR , \d[42]_BAR , \d[41]_BAR , \d[30] , 
        \d[22]_BAR , \d[46]_BAR , \d[35] , \d[19] , \d[10]_BAR , \d[8]_BAR , 
        \d[5]_BAR , \d[29] , \d[32] , \d[39]_BAR , \d[2] , \d[36]_BAR , 
        \d[25] , \d[13]_BAR , \d[38]_BAR , \d[20] , \d[18] , \d[17]_BAR , 
        \d[45]_BAR , \d[21] , \d[12] , \d[7] , \d[6] , \d[3]_BAR  );
  input [23:0] a;
  input [23:0] b;
  input clk, rst;
  output \d[47] , \d[44] , \d[43] , \d[40] , \d[37]_BAR , \d[34] , \d[31] ,
         \d[28] , \d[16] , \d[1] , \d[0] , \d[33]_BAR , \d[27]_BAR ,
         \d[26]_BAR , \d[24]_BAR , \d[23]_BAR , \d[15]_BAR , \d[14]_BAR ,
         \d[11]_BAR , \d[9]_BAR , \d[4]_BAR , \d[42]_BAR , \d[41]_BAR ,
         \d[30] , \d[22]_BAR , \d[46]_BAR , \d[35] , \d[19] , \d[10]_BAR ,
         \d[8]_BAR , \d[5]_BAR , \d[29] , \d[32] , \d[39]_BAR , \d[2] ,
         \d[36]_BAR , \d[25] , \d[13]_BAR , \d[38]_BAR , \d[20] , \d[18] ,
         \d[17]_BAR , \d[45]_BAR , \d[21] , \d[12] , \d[7] , \d[6] ,
         \d[3]_BAR ;
  wire   \intadd_0/A[4] , \intadd_0/A[3] , \intadd_0/A[2] , \intadd_0/A[1] ,
         \intadd_0/A[0] , \intadd_0/B[4] , \intadd_0/B[3] , \intadd_0/B[2] ,
         \intadd_0/B[1] , \intadd_0/B[0] , \intadd_0/CI , \intadd_0/SUM[2] ,
         \intadd_0/SUM[1] , \intadd_0/SUM[0] , \intadd_0/n5 , \intadd_0/n4 ,
         \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 , \intadd_1/A[4] ,
         \intadd_1/A[3] , \intadd_1/A[2] , \intadd_1/A[1] , \intadd_1/A[0] ,
         \intadd_1/B[4] , \intadd_1/B[3] , \intadd_1/B[2] , \intadd_1/B[1] ,
         \intadd_1/B[0] , \intadd_1/CI , \intadd_1/SUM[4] , \intadd_1/SUM[3] ,
         \intadd_1/SUM[2] , \intadd_1/SUM[1] , \intadd_1/SUM[0] ,
         \intadd_1/n5 , \intadd_1/n4 , \intadd_1/n3 , \intadd_1/n2 ,
         \intadd_1/n1 , \intadd_2/A[4] , \intadd_2/A[3] , \intadd_2/A[2] ,
         \intadd_2/A[1] , \intadd_2/A[0] , \intadd_2/B[4] , \intadd_2/B[3] ,
         \intadd_2/B[2] , \intadd_2/B[1] , \intadd_2/B[0] , \intadd_2/CI ,
         \intadd_2/SUM[4] , \intadd_2/SUM[2] , \intadd_2/SUM[0] ,
         \intadd_2/n5 , \intadd_2/n4 , \intadd_2/n3 , \intadd_2/n2 ,
         \intadd_2/n1 , \intadd_3/A[3] , \intadd_3/A[2] , \intadd_3/A[1] ,
         \intadd_3/A[0] , \intadd_3/B[1] , \intadd_3/B[0] , \intadd_3/CI ,
         \intadd_3/SUM[4] , \intadd_3/SUM[3] , \intadd_3/SUM[2] ,
         \intadd_3/SUM[1] , \intadd_3/SUM[0] , \intadd_3/n5 , \intadd_3/n4 ,
         \intadd_3/n3 , \intadd_3/n2 , \intadd_3/n1 , \intadd_4/A[1] ,
         \intadd_4/A[0] , \intadd_4/B[3] , \intadd_4/B[2] , \intadd_4/B[1] ,
         \intadd_4/B[0] , \intadd_4/CI , \intadd_4/SUM[4] , \intadd_4/SUM[3] ,
         \intadd_4/SUM[2] , \intadd_4/SUM[1] , \intadd_4/SUM[0] ,
         \intadd_4/n5 , \intadd_4/n4 , \intadd_4/n3 , \intadd_4/n2 ,
         \intadd_4/n1 , \intadd_5/A[4] , \intadd_5/A[3] , \intadd_5/A[2] ,
         \intadd_5/A[1] , \intadd_5/A[0] , \intadd_5/B[4] , \intadd_5/B[3] ,
         \intadd_5/B[2] , \intadd_5/B[1] , \intadd_5/B[0] , \intadd_5/CI ,
         \intadd_5/SUM[4] , \intadd_5/SUM[3] , \intadd_5/SUM[2] ,
         \intadd_5/SUM[1] , \intadd_5/SUM[0] , \intadd_5/n5 , \intadd_5/n4 ,
         \intadd_5/n3 , \intadd_5/n2 , \intadd_5/n1 , \intadd_6/A[4] ,
         \intadd_6/A[2] , \intadd_6/A[1] , \intadd_6/A[0] , \intadd_6/B[4] ,
         \intadd_6/B[3] , \intadd_6/B[2] , \intadd_6/B[1] , \intadd_6/B[0] ,
         \intadd_6/CI , \intadd_6/SUM[4] , \intadd_6/SUM[3] ,
         \intadd_6/SUM[2] , \intadd_6/SUM[1] , \intadd_6/SUM[0] ,
         \intadd_6/n5 , \intadd_6/n4 , \intadd_6/n3 , \intadd_6/n2 ,
         \intadd_6/n1 , \intadd_7/A[4] , \intadd_7/A[3] , \intadd_7/A[2] ,
         \intadd_7/A[1] , \intadd_7/A[0] , \intadd_7/B[3] , \intadd_7/B[2] ,
         \intadd_7/B[1] , \intadd_7/B[0] , \intadd_7/CI , \intadd_7/SUM[4] ,
         \intadd_7/SUM[3] , \intadd_7/SUM[2] , \intadd_7/SUM[1] ,
         \intadd_7/SUM[0] , \intadd_7/n5 , \intadd_7/n4 , \intadd_7/n3 ,
         \intadd_7/n2 , \intadd_7/n1 , \intadd_8/A[4] , \intadd_8/A[1] ,
         \intadd_8/A[0] , \intadd_8/B[4] , \intadd_8/B[1] , \intadd_8/B[0] ,
         \intadd_8/CI , \intadd_8/SUM[4] , \intadd_8/SUM[1] ,
         \intadd_8/SUM[0] , \intadd_8/n5 , \intadd_8/n4 , \intadd_8/n2 ,
         \intadd_8/n1 , \intadd_9/A[4] , \intadd_9/A[3] , \intadd_9/A[2] ,
         \intadd_9/A[1] , \intadd_9/A[0] , \intadd_9/B[4] , \intadd_9/B[3] ,
         \intadd_9/B[2] , \intadd_9/B[1] , \intadd_9/B[0] , \intadd_9/CI ,
         \intadd_9/SUM[4] , \intadd_9/SUM[3] , \intadd_9/SUM[2] ,
         \intadd_9/SUM[1] , \intadd_9/SUM[0] , \intadd_9/n5 , \intadd_9/n4 ,
         \intadd_9/n3 , \intadd_9/n2 , \intadd_9/n1 , \intadd_10/A[4] ,
         \intadd_10/A[3] , \intadd_10/A[2] , \intadd_10/A[1] ,
         \intadd_10/A[0] , \intadd_10/B[4] , \intadd_10/B[3] ,
         \intadd_10/B[2] , \intadd_10/B[1] , \intadd_10/B[0] , \intadd_10/CI ,
         \intadd_10/SUM[4] , \intadd_10/SUM[2] , \intadd_10/SUM[1] ,
         \intadd_10/n5 , \intadd_10/n4 , \intadd_10/n3 , \intadd_10/n2 ,
         \intadd_10/n1 , \intadd_11/A[1] , \intadd_11/B[3] , \intadd_11/B[0] ,
         \intadd_11/CI , \intadd_11/SUM[1] , \intadd_11/SUM[0] ,
         \intadd_11/n4 , \intadd_11/n3 , \intadd_11/n2 , \intadd_11/n1 ,
         \intadd_12/A[3] , \intadd_12/A[2] , \intadd_12/A[1] ,
         \intadd_12/A[0] , \intadd_12/B[3] , \intadd_12/B[2] ,
         \intadd_12/B[1] , \intadd_12/B[0] , \intadd_12/CI ,
         \intadd_12/SUM[3] , \intadd_12/SUM[2] , \intadd_12/SUM[1] ,
         \intadd_12/SUM[0] , \intadd_12/n4 , \intadd_12/n3 , \intadd_12/n2 ,
         \intadd_12/n1 , \intadd_13/A[3] , \intadd_13/A[2] , \intadd_13/A[1] ,
         \intadd_13/A[0] , \intadd_13/B[3] , \intadd_13/B[2] ,
         \intadd_13/B[1] , \intadd_13/B[0] , \intadd_13/CI ,
         \intadd_13/SUM[3] , \intadd_13/SUM[0] , \intadd_13/n4 ,
         \intadd_13/n3 , \intadd_13/n2 , \intadd_13/n1 , \intadd_14/A[3] ,
         \intadd_14/A[2] , \intadd_14/A[1] , \intadd_14/A[0] ,
         \intadd_14/B[3] , \intadd_14/B[2] , \intadd_14/B[1] ,
         \intadd_14/B[0] , \intadd_14/CI , \intadd_14/SUM[3] ,
         \intadd_14/SUM[0] , \intadd_14/n4 , \intadd_14/n3 , \intadd_14/n2 ,
         \intadd_14/n1 , \intadd_15/A[3] , \intadd_15/A[2] , \intadd_15/A[1] ,
         \intadd_15/A[0] , \intadd_15/B[3] , \intadd_15/B[2] ,
         \intadd_15/B[1] , \intadd_15/B[0] , \intadd_15/CI ,
         \intadd_15/SUM[0] , \intadd_15/n4 , \intadd_15/n3 , \intadd_15/n2 ,
         \intadd_15/n1 , \intadd_16/A[3] , \intadd_16/A[2] , \intadd_16/A[1] ,
         \intadd_16/A[0] , \intadd_16/B[3] , \intadd_16/B[2] ,
         \intadd_16/B[1] , \intadd_16/B[0] , \intadd_16/CI , \intadd_16/n4 ,
         \intadd_16/n3 , \intadd_16/n2 , \intadd_16/n1 , \intadd_17/A[1] ,
         \intadd_17/A[0] , \intadd_17/B[3] , \intadd_17/B[2] ,
         \intadd_17/B[1] , \intadd_17/B[0] , \intadd_17/CI ,
         \intadd_17/SUM[3] , \intadd_17/SUM[1] , \intadd_17/SUM[0] ,
         \intadd_17/n4 , \intadd_17/n3 , \intadd_17/n2 , \intadd_17/n1 ,
         \intadd_18/A[3] , \intadd_18/A[2] , \intadd_18/A[1] ,
         \intadd_18/A[0] , \intadd_18/B[3] , \intadd_18/B[2] ,
         \intadd_18/B[1] , \intadd_18/B[0] , \intadd_18/CI ,
         \intadd_18/SUM[2] , \intadd_18/n4 , \intadd_18/n3 , \intadd_18/n2 ,
         \intadd_18/n1 , \intadd_19/A[3] , \intadd_19/A[2] , \intadd_19/A[1] ,
         \intadd_19/A[0] , \intadd_19/B[3] , \intadd_19/B[2] ,
         \intadd_19/B[1] , \intadd_19/B[0] , \intadd_19/CI ,
         \intadd_19/SUM[3] , \intadd_19/SUM[2] , \intadd_19/SUM[1] ,
         \intadd_19/SUM[0] , \intadd_19/n4 , \intadd_19/n3 , \intadd_19/n2 ,
         \intadd_19/n1 , \intadd_20/A[3] , \intadd_20/A[2] , \intadd_20/A[1] ,
         \intadd_20/A[0] , \intadd_20/B[2] , \intadd_20/B[1] ,
         \intadd_20/B[0] , \intadd_20/CI , \intadd_20/SUM[3] ,
         \intadd_20/SUM[2] , \intadd_20/n4 , \intadd_20/n3 , \intadd_20/n2 ,
         \intadd_20/n1 , \intadd_21/A[3] , \intadd_21/A[2] , \intadd_21/A[1] ,
         \intadd_21/A[0] , \intadd_21/B[2] , \intadd_21/B[1] ,
         \intadd_21/B[0] , \intadd_21/CI , \intadd_21/SUM[3] ,
         \intadd_21/SUM[2] , \intadd_21/SUM[1] , \intadd_21/SUM[0] ,
         \intadd_21/n4 , \intadd_21/n3 , \intadd_21/n2 , \intadd_21/n1 ,
         \intadd_22/A[3] , \intadd_22/A[2] , \intadd_22/A[1] ,
         \intadd_22/A[0] , \intadd_22/B[3] , \intadd_22/B[2] ,
         \intadd_22/B[1] , \intadd_22/B[0] , \intadd_22/CI ,
         \intadd_22/SUM[3] , \intadd_22/SUM[2] , \intadd_22/SUM[1] ,
         \intadd_22/SUM[0] , \intadd_22/n4 , \intadd_22/n3 , \intadd_22/n2 ,
         \intadd_22/n1 , \intadd_23/A[3] , \intadd_23/A[2] , \intadd_23/A[1] ,
         \intadd_23/A[0] , \intadd_23/B[2] , \intadd_23/B[1] ,
         \intadd_23/B[0] , \intadd_23/CI , \intadd_23/SUM[3] ,
         \intadd_23/SUM[2] , \intadd_23/SUM[1] , \intadd_23/SUM[0] ,
         \intadd_23/n4 , \intadd_23/n3 , \intadd_23/n2 , \intadd_23/n1 ,
         \intadd_24/A[2] , \intadd_24/A[1] , \intadd_24/A[0] ,
         \intadd_24/B[2] , \intadd_24/B[1] , \intadd_24/B[0] , \intadd_24/CI ,
         \intadd_24/n3 , \intadd_24/n2 , \intadd_24/n1 , \intadd_25/A[1] ,
         \intadd_25/A[0] , \intadd_25/B[2] , \intadd_25/B[1] ,
         \intadd_25/B[0] , \intadd_25/CI , \intadd_25/SUM[2] ,
         \intadd_25/SUM[1] , \intadd_25/SUM[0] , \intadd_25/n3 ,
         \intadd_25/n2 , \intadd_25/n1 , \intadd_26/A[2] , \intadd_26/A[1] ,
         \intadd_26/A[0] , \intadd_26/B[2] , \intadd_26/B[1] ,
         \intadd_26/B[0] , \intadd_26/CI , \intadd_26/SUM[2] ,
         \intadd_26/SUM[1] , \intadd_26/SUM[0] , \intadd_26/n3 ,
         \intadd_26/n2 , \intadd_26/n1 , \intadd_27/A[1] , \intadd_27/A[0] ,
         \intadd_27/B[2] , \intadd_27/B[1] , \intadd_27/B[0] , \intadd_27/CI ,
         \intadd_27/SUM[1] , \intadd_27/SUM[0] , \intadd_27/n3 ,
         \intadd_27/n2 , \intadd_27/n1 , \intadd_28/A[2] , \intadd_28/A[1] ,
         \intadd_28/A[0] , \intadd_28/B[2] , \intadd_28/B[1] ,
         \intadd_28/B[0] , \intadd_28/CI , \intadd_28/SUM[2] ,
         \intadd_28/SUM[1] , \intadd_28/SUM[0] , \intadd_28/n3 ,
         \intadd_28/n2 , \intadd_28/n1 , \intadd_29/A[2] , \intadd_29/A[1] ,
         \intadd_29/A[0] , \intadd_29/B[1] , \intadd_29/B[0] , \intadd_29/CI ,
         \intadd_29/SUM[1] , \intadd_29/SUM[0] , \intadd_29/n3 ,
         \intadd_29/n2 , \intadd_29/n1 , \intadd_30/A[2] , \intadd_30/A[1] ,
         \intadd_30/A[0] , \intadd_30/B[2] , \intadd_30/B[1] ,
         \intadd_30/B[0] , \intadd_30/CI , \intadd_30/SUM[2] ,
         \intadd_30/SUM[1] , \intadd_30/SUM[0] , \intadd_30/n3 ,
         \intadd_30/n2 , \intadd_30/n1 , \intadd_31/A[1] , \intadd_31/A[0] ,
         \intadd_31/B[0] , \intadd_31/SUM[2] , \intadd_31/SUM[1] ,
         \intadd_31/n3 , \intadd_31/n2 , \intadd_31/n1 , \intadd_32/A[2] ,
         \intadd_32/A[1] , \intadd_32/A[0] , \intadd_32/B[2] ,
         \intadd_32/B[1] , \intadd_32/B[0] , \intadd_32/CI ,
         \intadd_32/SUM[2] , \intadd_32/SUM[1] , \intadd_32/SUM[0] ,
         \intadd_32/n3 , \intadd_32/n2 , \intadd_32/n1 , \intadd_33/A[2] ,
         \intadd_33/A[0] , \intadd_33/B[2] , \intadd_33/B[1] ,
         \intadd_33/B[0] , \intadd_33/CI , \intadd_33/SUM[0] , \intadd_33/n3 ,
         \intadd_33/n2 , \intadd_33/n1 , \intadd_34/A[2] , \intadd_34/A[1] ,
         \intadd_34/A[0] , \intadd_34/B[2] , \intadd_34/B[1] ,
         \intadd_34/B[0] , \intadd_34/CI , \intadd_34/n3 , \intadd_34/n2 ,
         \intadd_34/n1 , \intadd_35/A[0] , \intadd_35/B[2] , \intadd_35/B[1] ,
         \intadd_35/B[0] , \intadd_35/CI , \intadd_35/SUM[2] ,
         \intadd_35/SUM[0] , \intadd_35/n3 , \intadd_35/n2 , \intadd_35/n1 ,
         n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281;
  assign \d[12]  = \intadd_8/SUM[4] ;
  assign \d[45]_BAR  = \intadd_12/SUM[3] ;
  assign \d[7]  = \intadd_26/SUM[2] ;
  assign \d[6]  = \intadd_26/SUM[1] ;

  FA_X1 \intadd_0/U6  ( .A(\intadd_0/A[0] ), .B(\intadd_0/B[0] ), .CI(
        \intadd_0/CI ), .CO(\intadd_0/n5 ), .S(\intadd_0/SUM[0] ) );
  FA_X1 \intadd_0/U5  ( .A(\intadd_0/A[1] ), .B(\intadd_0/B[1] ), .CI(
        \intadd_0/n5 ), .CO(\intadd_0/n4 ), .S(\intadd_0/SUM[1] ) );
  FA_X1 \intadd_0/U4  ( .A(\intadd_0/A[2] ), .B(\intadd_0/B[2] ), .CI(
        \intadd_0/n4 ), .CO(\intadd_0/n3 ), .S(\intadd_0/SUM[2] ) );
  FA_X1 \intadd_0/U3  ( .A(\intadd_0/A[3] ), .B(\intadd_0/B[3] ), .CI(
        \intadd_0/n3 ), .CO(\intadd_0/n2 ), .S(\d[13]_BAR ) );
  FA_X1 \intadd_0/U2  ( .A(\intadd_0/A[4] ), .B(\intadd_0/B[4] ), .CI(
        \intadd_0/n2 ), .CO(\intadd_0/n1 ), .S(\d[14]_BAR ) );
  FA_X1 \intadd_1/U6  ( .A(\intadd_1/A[0] ), .B(\intadd_1/B[0] ), .CI(
        \intadd_1/CI ), .CO(\intadd_1/n5 ), .S(\intadd_1/SUM[0] ) );
  FA_X1 \intadd_1/U5  ( .A(\intadd_1/A[1] ), .B(\intadd_1/B[1] ), .CI(
        \intadd_1/n5 ), .CO(\intadd_1/n4 ), .S(\intadd_1/SUM[1] ) );
  FA_X1 \intadd_1/U4  ( .A(\intadd_1/A[2] ), .B(\intadd_1/B[2] ), .CI(
        \intadd_1/n4 ), .CO(\intadd_1/n3 ), .S(\intadd_1/SUM[2] ) );
  FA_X1 \intadd_1/U3  ( .A(\intadd_1/A[3] ), .B(\intadd_1/B[3] ), .CI(
        \intadd_1/n3 ), .CO(\intadd_1/n2 ), .S(\intadd_1/SUM[3] ) );
  FA_X1 \intadd_1/U2  ( .A(\intadd_1/A[4] ), .B(\intadd_1/B[4] ), .CI(
        \intadd_1/n2 ), .CO(\intadd_1/n1 ), .S(\intadd_1/SUM[4] ) );
  FA_X1 \intadd_2/U6  ( .A(\intadd_2/A[0] ), .B(\intadd_2/B[0] ), .CI(
        \intadd_2/CI ), .CO(\intadd_2/n5 ), .S(\intadd_2/SUM[0] ) );
  FA_X1 \intadd_2/U5  ( .A(\intadd_2/A[1] ), .B(\intadd_2/B[1] ), .CI(
        \intadd_2/n5 ), .CO(\intadd_2/n4 ), .S(\intadd_1/A[2] ) );
  FA_X1 \intadd_2/U4  ( .A(\intadd_2/A[2] ), .B(\intadd_2/B[2] ), .CI(
        \intadd_2/n4 ), .CO(\intadd_2/n3 ), .S(\intadd_2/SUM[2] ) );
  FA_X1 \intadd_2/U3  ( .A(\intadd_2/A[3] ), .B(\intadd_2/B[3] ), .CI(
        \intadd_2/n3 ), .CO(\intadd_2/n2 ), .S(\intadd_1/A[4] ) );
  FA_X1 \intadd_2/U2  ( .A(\intadd_2/A[4] ), .B(\intadd_2/B[4] ), .CI(
        \intadd_2/n2 ), .CO(\intadd_2/n1 ), .S(\intadd_2/SUM[4] ) );
  FA_X1 \intadd_3/U6  ( .A(\intadd_3/A[0] ), .B(\intadd_3/B[0] ), .CI(
        \intadd_3/CI ), .CO(\intadd_3/n5 ), .S(\intadd_3/SUM[0] ) );
  FA_X1 \intadd_3/U5  ( .A(\intadd_3/A[1] ), .B(\intadd_3/B[1] ), .CI(
        \intadd_3/n5 ), .CO(\intadd_3/n4 ), .S(\intadd_3/SUM[1] ) );
  FA_X1 \intadd_3/U4  ( .A(\intadd_3/A[2] ), .B(\intadd_2/SUM[0] ), .CI(
        \intadd_3/n4 ), .CO(\intadd_3/n3 ), .S(\intadd_3/SUM[2] ) );
  FA_X1 \intadd_3/U3  ( .A(\intadd_3/A[3] ), .B(\intadd_25/n1 ), .CI(
        \intadd_3/n3 ), .CO(\intadd_3/n2 ), .S(\intadd_3/SUM[3] ) );
  FA_X1 \intadd_3/U2  ( .A(\intadd_1/SUM[3] ), .B(\intadd_2/SUM[2] ), .CI(
        \intadd_3/n2 ), .CO(\intadd_3/n1 ), .S(\intadd_3/SUM[4] ) );
  FA_X1 \intadd_4/U6  ( .A(\intadd_4/A[0] ), .B(\intadd_4/B[0] ), .CI(
        \intadd_4/CI ), .CO(\intadd_4/n5 ), .S(\intadd_4/SUM[0] ) );
  FA_X1 \intadd_4/U5  ( .A(\intadd_4/A[1] ), .B(\intadd_4/B[1] ), .CI(
        \intadd_4/n5 ), .CO(\intadd_4/n4 ), .S(\intadd_4/SUM[1] ) );
  FA_X1 \intadd_4/U4  ( .A(\intadd_1/SUM[0] ), .B(\intadd_4/B[2] ), .CI(
        \intadd_4/n4 ), .CO(\intadd_4/n3 ), .S(\intadd_4/SUM[2] ) );
  FA_X1 \intadd_4/U3  ( .A(\intadd_3/SUM[2] ), .B(\intadd_4/B[3] ), .CI(
        \intadd_4/n3 ), .CO(\intadd_4/n2 ), .S(\intadd_4/SUM[3] ) );
  FA_X1 \intadd_4/U2  ( .A(\intadd_1/SUM[2] ), .B(\intadd_3/SUM[3] ), .CI(
        \intadd_4/n2 ), .CO(\intadd_4/n1 ), .S(\intadd_4/SUM[4] ) );
  FA_X1 \intadd_5/U6  ( .A(\intadd_5/A[0] ), .B(\intadd_5/B[0] ), .CI(
        \intadd_5/CI ), .CO(\intadd_5/n5 ), .S(\intadd_5/SUM[0] ) );
  FA_X1 \intadd_5/U5  ( .A(\intadd_5/A[1] ), .B(\intadd_5/B[1] ), .CI(
        \intadd_5/n5 ), .CO(\intadd_5/n4 ), .S(\intadd_5/SUM[1] ) );
  FA_X1 \intadd_5/U4  ( .A(\intadd_5/A[2] ), .B(\intadd_5/B[2] ), .CI(
        \intadd_5/n4 ), .CO(\intadd_5/n3 ), .S(\intadd_5/SUM[2] ) );
  FA_X1 \intadd_5/U3  ( .A(\intadd_5/A[3] ), .B(\intadd_5/B[3] ), .CI(
        \intadd_5/n3 ), .CO(\intadd_5/n2 ), .S(\intadd_5/SUM[3] ) );
  FA_X1 \intadd_5/U2  ( .A(\intadd_5/A[4] ), .B(\intadd_5/B[4] ), .CI(
        \intadd_5/n2 ), .CO(\intadd_5/n1 ), .S(\intadd_5/SUM[4] ) );
  FA_X1 \intadd_6/U6  ( .A(\intadd_6/A[0] ), .B(\intadd_6/B[0] ), .CI(
        \intadd_6/CI ), .CO(\intadd_6/n5 ), .S(\intadd_6/SUM[0] ) );
  FA_X1 \intadd_6/U5  ( .A(\intadd_6/A[1] ), .B(\intadd_6/B[1] ), .CI(
        \intadd_6/n5 ), .CO(\intadd_6/n4 ), .S(\intadd_6/SUM[1] ) );
  FA_X1 \intadd_6/U4  ( .A(\intadd_6/A[2] ), .B(\intadd_6/B[2] ), .CI(
        \intadd_6/n4 ), .CO(\intadd_6/n3 ), .S(\intadd_6/SUM[2] ) );
  FA_X1 \intadd_6/U3  ( .A(\intadd_24/n1 ), .B(\intadd_6/B[3] ), .CI(
        \intadd_6/n3 ), .CO(\intadd_6/n2 ), .S(\intadd_6/SUM[3] ) );
  FA_X1 \intadd_6/U2  ( .A(\intadd_6/A[4] ), .B(\intadd_6/B[4] ), .CI(
        \intadd_6/n2 ), .CO(\intadd_6/n1 ), .S(\intadd_6/SUM[4] ) );
  FA_X1 \intadd_7/U6  ( .A(\intadd_7/A[0] ), .B(\intadd_7/B[0] ), .CI(
        \intadd_7/CI ), .CO(\intadd_7/n5 ), .S(\intadd_7/SUM[0] ) );
  FA_X1 \intadd_7/U5  ( .A(\intadd_7/A[1] ), .B(\intadd_7/B[1] ), .CI(
        \intadd_7/n5 ), .CO(\intadd_7/n4 ), .S(\intadd_7/SUM[1] ) );
  FA_X1 \intadd_7/U4  ( .A(\intadd_7/A[2] ), .B(\intadd_7/B[2] ), .CI(
        \intadd_7/n4 ), .CO(\intadd_7/n3 ), .S(\intadd_7/SUM[2] ) );
  FA_X1 \intadd_7/U3  ( .A(\intadd_7/A[3] ), .B(\intadd_7/B[3] ), .CI(
        \intadd_7/n3 ), .CO(\intadd_7/n2 ), .S(\intadd_7/SUM[3] ) );
  FA_X1 \intadd_7/U2  ( .A(\intadd_7/A[4] ), .B(\intadd_6/SUM[3] ), .CI(
        \intadd_7/n2 ), .CO(\intadd_7/n1 ), .S(\intadd_7/SUM[4] ) );
  FA_X1 \intadd_8/U6  ( .A(\intadd_8/A[0] ), .B(\intadd_8/B[0] ), .CI(
        \intadd_8/CI ), .CO(\intadd_8/n5 ), .S(\intadd_8/SUM[0] ) );
  FA_X1 \intadd_8/U5  ( .A(\intadd_8/A[1] ), .B(\intadd_8/B[1] ), .CI(
        \intadd_8/n5 ), .CO(\intadd_8/n4 ), .S(\intadd_8/SUM[1] ) );
  FA_X1 \intadd_8/U2  ( .A(\intadd_8/A[4] ), .B(\intadd_8/B[4] ), .CI(
        \intadd_8/n2 ), .CO(\intadd_8/n1 ), .S(\intadd_8/SUM[4] ) );
  FA_X1 \intadd_9/U6  ( .A(\intadd_9/A[0] ), .B(\intadd_9/B[0] ), .CI(
        \intadd_9/CI ), .CO(\intadd_9/n5 ), .S(\intadd_9/SUM[0] ) );
  FA_X1 \intadd_9/U5  ( .A(\intadd_9/A[1] ), .B(\intadd_9/B[1] ), .CI(
        \intadd_9/n5 ), .CO(\intadd_9/n4 ), .S(\intadd_9/SUM[1] ) );
  FA_X1 \intadd_9/U4  ( .A(\intadd_9/A[2] ), .B(\intadd_9/B[2] ), .CI(
        \intadd_9/n4 ), .CO(\intadd_9/n3 ), .S(\intadd_9/SUM[2] ) );
  FA_X1 \intadd_9/U3  ( .A(\intadd_9/A[3] ), .B(\intadd_9/B[3] ), .CI(
        \intadd_9/n3 ), .CO(\intadd_9/n2 ), .S(\intadd_9/SUM[3] ) );
  FA_X1 \intadd_9/U2  ( .A(\intadd_9/A[4] ), .B(\intadd_9/B[4] ), .CI(
        \intadd_9/n2 ), .CO(\intadd_9/n1 ), .S(\intadd_9/SUM[4] ) );
  FA_X1 \intadd_10/U6  ( .A(\intadd_10/A[0] ), .B(\intadd_10/B[0] ), .CI(
        \intadd_10/CI ), .CO(\intadd_10/n5 ), .S(\intadd_9/A[1] ) );
  FA_X1 \intadd_10/U5  ( .A(\intadd_10/A[1] ), .B(\intadd_10/B[1] ), .CI(
        \intadd_10/n5 ), .CO(\intadd_10/n4 ), .S(\intadd_10/SUM[1] ) );
  FA_X1 \intadd_10/U4  ( .A(\intadd_10/A[2] ), .B(\intadd_10/B[2] ), .CI(
        \intadd_10/n4 ), .CO(\intadd_10/n3 ), .S(\intadd_10/SUM[2] ) );
  FA_X1 \intadd_10/U3  ( .A(\intadd_10/A[3] ), .B(\intadd_10/B[3] ), .CI(
        \intadd_10/n3 ), .CO(\intadd_10/n2 ), .S(\intadd_9/A[4] ) );
  FA_X1 \intadd_10/U2  ( .A(\intadd_10/A[4] ), .B(\intadd_10/B[4] ), .CI(
        \intadd_10/n2 ), .CO(\intadd_10/n1 ), .S(\intadd_10/SUM[4] ) );
  FA_X1 \intadd_11/U5  ( .A(\intadd_31/n1 ), .B(\intadd_11/B[0] ), .CI(
        \intadd_11/CI ), .CO(\intadd_11/n4 ), .S(\intadd_11/SUM[0] ) );
  FA_X1 \intadd_11/U4  ( .A(\intadd_11/A[1] ), .B(\intadd_9/SUM[4] ), .CI(
        \intadd_11/n4 ), .CO(\intadd_11/n3 ), .S(\intadd_11/SUM[1] ) );
  FA_X1 \intadd_11/U3  ( .A(\intadd_9/n1 ), .B(\intadd_10/SUM[4] ), .CI(
        \intadd_11/n3 ), .CO(\intadd_11/n2 ), .S(\d[22]_BAR ) );
  FA_X1 \intadd_11/U2  ( .A(\intadd_10/n1 ), .B(\intadd_11/B[3] ), .CI(
        \intadd_11/n2 ), .CO(\intadd_11/n1 ), .S(\d[23]_BAR ) );
  FA_X1 \intadd_12/U5  ( .A(\intadd_12/A[0] ), .B(\intadd_12/B[0] ), .CI(
        \intadd_12/CI ), .CO(\intadd_12/n4 ), .S(\intadd_12/SUM[0] ) );
  FA_X1 \intadd_12/U4  ( .A(\intadd_12/A[1] ), .B(\intadd_12/B[1] ), .CI(
        \intadd_12/n4 ), .CO(\intadd_12/n3 ), .S(\intadd_12/SUM[1] ) );
  FA_X1 \intadd_12/U3  ( .A(\intadd_12/A[2] ), .B(\intadd_12/B[2] ), .CI(
        \intadd_12/n3 ), .CO(\intadd_12/n2 ), .S(\intadd_12/SUM[2] ) );
  FA_X1 \intadd_12/U2  ( .A(\intadd_12/A[3] ), .B(\intadd_12/n2 ), .CI(
        \intadd_12/B[3] ), .CO(\intadd_12/n1 ), .S(\intadd_12/SUM[3] ) );
  FA_X1 \intadd_13/U5  ( .A(\intadd_13/A[0] ), .B(\intadd_13/B[0] ), .CI(
        \intadd_13/CI ), .CO(\intadd_13/n4 ), .S(\intadd_13/SUM[0] ) );
  FA_X1 \intadd_13/U4  ( .A(\intadd_13/A[1] ), .B(\intadd_13/B[1] ), .CI(
        \intadd_13/n4 ), .CO(\intadd_13/n3 ), .S(\intadd_2/A[3] ) );
  FA_X1 \intadd_13/U3  ( .A(\intadd_13/A[2] ), .B(\intadd_13/B[2] ), .CI(
        \intadd_13/n3 ), .CO(\intadd_13/n2 ), .S(\intadd_2/A[4] ) );
  FA_X1 \intadd_13/U2  ( .A(\intadd_13/A[3] ), .B(\intadd_13/B[3] ), .CI(
        \intadd_13/n2 ), .CO(\intadd_13/n1 ), .S(\intadd_13/SUM[3] ) );
  FA_X1 \intadd_14/U5  ( .A(\intadd_14/A[0] ), .B(\intadd_14/B[0] ), .CI(
        \intadd_14/CI ), .CO(\intadd_14/n4 ), .S(\intadd_14/SUM[0] ) );
  FA_X1 \intadd_14/U4  ( .A(\intadd_14/A[1] ), .B(\intadd_14/B[1] ), .CI(
        \intadd_14/n4 ), .CO(\intadd_14/n3 ), .S(\intadd_13/B[2] ) );
  FA_X1 \intadd_14/U3  ( .A(\intadd_14/A[2] ), .B(\intadd_14/B[2] ), .CI(
        \intadd_14/n3 ), .CO(\intadd_14/n2 ), .S(\intadd_13/A[3] ) );
  FA_X1 \intadd_14/U2  ( .A(\intadd_14/A[3] ), .B(\intadd_14/B[3] ), .CI(
        \intadd_14/n2 ), .CO(\intadd_14/n1 ), .S(\intadd_14/SUM[3] ) );
  FA_X1 \intadd_15/U5  ( .A(\intadd_15/A[0] ), .B(\intadd_15/B[0] ), .CI(
        \intadd_15/CI ), .CO(\intadd_15/n4 ), .S(\intadd_15/SUM[0] ) );
  FA_X1 \intadd_15/U4  ( .A(\intadd_15/A[1] ), .B(\intadd_15/B[1] ), .CI(
        \intadd_15/n4 ), .CO(\intadd_15/n3 ), .S(\intadd_5/A[2] ) );
  FA_X1 \intadd_15/U3  ( .A(\intadd_15/A[2] ), .B(\intadd_15/B[2] ), .CI(
        \intadd_15/n3 ), .CO(\intadd_15/n2 ), .S(\intadd_5/A[3] ) );
  FA_X1 \intadd_15/U2  ( .A(\intadd_15/A[3] ), .B(\intadd_15/B[3] ), .CI(
        \intadd_15/n2 ), .CO(\intadd_15/n1 ), .S(\intadd_5/A[4] ) );
  FA_X1 \intadd_16/U5  ( .A(\intadd_16/A[0] ), .B(\intadd_16/B[0] ), .CI(
        \intadd_16/CI ), .CO(\intadd_16/n4 ), .S(\intadd_6/A[1] ) );
  FA_X1 \intadd_16/U4  ( .A(\intadd_16/A[1] ), .B(\intadd_16/B[1] ), .CI(
        \intadd_16/n4 ), .CO(\intadd_16/n3 ), .S(\intadd_6/B[2] ) );
  FA_X1 \intadd_16/U3  ( .A(\intadd_16/A[2] ), .B(\intadd_16/B[2] ), .CI(
        \intadd_16/n3 ), .CO(\intadd_16/n2 ), .S(\intadd_6/B[3] ) );
  FA_X1 \intadd_16/U2  ( .A(\intadd_16/A[3] ), .B(\intadd_16/B[3] ), .CI(
        \intadd_16/n2 ), .CO(\intadd_16/n1 ), .S(\intadd_6/B[4] ) );
  FA_X1 \intadd_17/U5  ( .A(\intadd_17/A[0] ), .B(\intadd_17/B[0] ), .CI(
        \intadd_17/CI ), .CO(\intadd_17/n4 ), .S(\intadd_17/SUM[0] ) );
  FA_X1 \intadd_17/U4  ( .A(\intadd_17/A[1] ), .B(\intadd_17/B[1] ), .CI(
        \intadd_17/n4 ), .CO(\intadd_17/n3 ), .S(\intadd_17/SUM[1] ) );
  FA_X1 \intadd_17/U3  ( .A(\intadd_3/SUM[0] ), .B(\intadd_17/B[2] ), .CI(
        \intadd_17/n3 ), .CO(\intadd_17/n2 ), .S(\intadd_15/A[3] ) );
  FA_X1 \intadd_17/U2  ( .A(\intadd_4/SUM[2] ), .B(\intadd_17/B[3] ), .CI(
        \intadd_17/n2 ), .CO(\intadd_17/n1 ), .S(\intadd_17/SUM[3] ) );
  FA_X1 \intadd_18/U5  ( .A(\intadd_18/A[0] ), .B(\intadd_18/B[0] ), .CI(
        \intadd_18/CI ), .CO(\intadd_18/n4 ), .S(\intadd_0/B[1] ) );
  FA_X1 \intadd_18/U4  ( .A(\intadd_18/A[1] ), .B(\intadd_18/B[1] ), .CI(
        \intadd_18/n4 ), .CO(\intadd_18/n3 ), .S(\intadd_0/B[2] ) );
  FA_X1 \intadd_18/U3  ( .A(\intadd_18/A[2] ), .B(\intadd_18/B[2] ), .CI(
        \intadd_18/n3 ), .CO(\intadd_18/n2 ), .S(\intadd_18/SUM[2] ) );
  FA_X1 \intadd_18/U2  ( .A(\intadd_18/A[3] ), .B(\intadd_18/B[3] ), .CI(
        \intadd_18/n2 ), .CO(\intadd_18/n1 ), .S(\intadd_0/A[4] ) );
  FA_X1 \intadd_19/U5  ( .A(\intadd_19/A[0] ), .B(\intadd_19/B[0] ), .CI(
        \intadd_19/CI ), .CO(\intadd_19/n4 ), .S(\intadd_19/SUM[0] ) );
  FA_X1 \intadd_19/U4  ( .A(\intadd_19/A[1] ), .B(\intadd_19/B[1] ), .CI(
        \intadd_19/n4 ), .CO(\intadd_19/n3 ), .S(\intadd_19/SUM[1] ) );
  FA_X1 \intadd_19/U3  ( .A(\intadd_19/A[2] ), .B(\intadd_19/B[2] ), .CI(
        \intadd_19/n3 ), .CO(\intadd_19/n2 ), .S(\intadd_19/SUM[2] ) );
  FA_X1 \intadd_19/U2  ( .A(\intadd_19/A[3] ), .B(\intadd_19/B[3] ), .CI(
        \intadd_19/n2 ), .CO(\intadd_19/n1 ), .S(\intadd_19/SUM[3] ) );
  FA_X1 \intadd_20/U5  ( .A(\intadd_20/A[0] ), .B(\intadd_20/B[0] ), .CI(
        \intadd_20/CI ), .CO(\intadd_20/n4 ), .S(\intadd_18/B[2] ) );
  FA_X1 \intadd_20/U4  ( .A(\intadd_20/A[1] ), .B(\intadd_20/B[1] ), .CI(
        \intadd_20/n4 ), .CO(\intadd_20/n3 ), .S(\intadd_18/A[3] ) );
  FA_X1 \intadd_20/U3  ( .A(\intadd_20/A[2] ), .B(\intadd_20/B[2] ), .CI(
        \intadd_20/n3 ), .CO(\intadd_20/n2 ), .S(\intadd_20/SUM[2] ) );
  FA_X1 \intadd_20/U2  ( .A(\intadd_20/A[3] ), .B(\intadd_19/SUM[2] ), .CI(
        \intadd_20/n2 ), .CO(\intadd_20/n1 ), .S(\intadd_20/SUM[3] ) );
  FA_X1 \intadd_21/U5  ( .A(\intadd_21/A[0] ), .B(\intadd_21/B[0] ), .CI(
        \intadd_21/CI ), .CO(\intadd_21/n4 ), .S(\intadd_21/SUM[0] ) );
  FA_X1 \intadd_21/U4  ( .A(\intadd_21/A[1] ), .B(\intadd_21/B[1] ), .CI(
        \intadd_21/n4 ), .CO(\intadd_21/n3 ), .S(\intadd_21/SUM[1] ) );
  FA_X1 \intadd_21/U3  ( .A(\intadd_21/A[2] ), .B(\intadd_21/B[2] ), .CI(
        \intadd_21/n3 ), .CO(\intadd_21/n2 ), .S(\intadd_21/SUM[2] ) );
  FA_X1 \intadd_21/U2  ( .A(\intadd_21/A[3] ), .B(\intadd_10/SUM[1] ), .CI(
        \intadd_21/n2 ), .CO(\intadd_21/n1 ), .S(\intadd_21/SUM[3] ) );
  FA_X1 \intadd_22/U5  ( .A(\intadd_22/A[0] ), .B(\intadd_22/B[0] ), .CI(
        \intadd_22/CI ), .CO(\intadd_22/n4 ), .S(\intadd_22/SUM[0] ) );
  FA_X1 \intadd_22/U4  ( .A(\intadd_22/A[1] ), .B(\intadd_22/B[1] ), .CI(
        \intadd_22/n4 ), .CO(\intadd_22/n3 ), .S(\intadd_22/SUM[1] ) );
  FA_X1 \intadd_22/U3  ( .A(\intadd_22/A[2] ), .B(\intadd_22/B[2] ), .CI(
        \intadd_22/n3 ), .CO(\intadd_22/n2 ), .S(\intadd_22/SUM[2] ) );
  FA_X1 \intadd_22/U2  ( .A(\intadd_22/A[3] ), .B(\intadd_22/B[3] ), .CI(
        \intadd_22/n2 ), .CO(\intadd_22/n1 ), .S(\intadd_22/SUM[3] ) );
  FA_X1 \intadd_23/U5  ( .A(\intadd_23/A[0] ), .B(\intadd_23/B[0] ), .CI(
        \intadd_23/CI ), .CO(\intadd_23/n4 ), .S(\intadd_23/SUM[0] ) );
  FA_X1 \intadd_23/U4  ( .A(\intadd_23/A[1] ), .B(\intadd_23/B[1] ), .CI(
        \intadd_23/n4 ), .CO(\intadd_23/n3 ), .S(\intadd_23/SUM[1] ) );
  FA_X1 \intadd_23/U3  ( .A(\intadd_23/A[2] ), .B(\intadd_23/B[2] ), .CI(
        \intadd_23/n3 ), .CO(\intadd_23/n2 ), .S(\intadd_23/SUM[2] ) );
  FA_X1 \intadd_23/U2  ( .A(\intadd_23/A[3] ), .B(\intadd_22/SUM[2] ), .CI(
        \intadd_23/n2 ), .CO(\intadd_23/n1 ), .S(\intadd_23/SUM[3] ) );
  FA_X1 \intadd_24/U4  ( .A(\intadd_24/A[0] ), .B(\intadd_24/B[0] ), .CI(
        \intadd_24/CI ), .CO(\intadd_24/n3 ), .S(\intadd_7/B[1] ) );
  FA_X1 \intadd_24/U3  ( .A(\intadd_24/A[1] ), .B(\intadd_24/B[1] ), .CI(
        \intadd_24/n3 ), .CO(\intadd_24/n2 ), .S(\intadd_7/B[2] ) );
  FA_X1 \intadd_24/U2  ( .A(\intadd_24/A[2] ), .B(\intadd_24/B[2] ), .CI(
        \intadd_24/n2 ), .CO(\intadd_24/n1 ), .S(\intadd_7/B[3] ) );
  FA_X1 \intadd_25/U4  ( .A(\intadd_25/A[0] ), .B(\intadd_25/B[0] ), .CI(
        \intadd_25/CI ), .CO(\intadd_25/n3 ), .S(\intadd_25/SUM[0] ) );
  FA_X1 \intadd_25/U3  ( .A(\intadd_25/A[1] ), .B(\intadd_25/B[1] ), .CI(
        \intadd_25/n3 ), .CO(\intadd_25/n2 ), .S(\intadd_25/SUM[1] ) );
  FA_X1 \intadd_25/U2  ( .A(\intadd_1/SUM[1] ), .B(\intadd_25/B[2] ), .CI(
        \intadd_25/n2 ), .CO(\intadd_25/n1 ), .S(\intadd_25/SUM[2] ) );
  FA_X1 \intadd_26/U4  ( .A(\intadd_26/A[0] ), .B(\intadd_26/B[0] ), .CI(
        \intadd_26/CI ), .CO(\intadd_26/n3 ), .S(\intadd_26/SUM[0] ) );
  FA_X1 \intadd_26/U3  ( .A(\intadd_26/A[1] ), .B(\intadd_26/B[1] ), .CI(
        \intadd_26/n3 ), .CO(\intadd_26/n2 ), .S(\intadd_26/SUM[1] ) );
  FA_X1 \intadd_26/U2  ( .A(\intadd_26/A[2] ), .B(\intadd_26/B[2] ), .CI(
        \intadd_26/n2 ), .CO(\intadd_26/n1 ), .S(\intadd_26/SUM[2] ) );
  FA_X1 \intadd_27/U4  ( .A(\intadd_27/A[0] ), .B(\intadd_27/B[0] ), .CI(
        \intadd_27/CI ), .CO(\intadd_27/n3 ), .S(\intadd_27/SUM[0] ) );
  FA_X1 \intadd_27/U3  ( .A(\intadd_27/A[1] ), .B(\intadd_27/B[1] ), .CI(
        \intadd_27/n3 ), .CO(\intadd_27/n2 ), .S(\intadd_27/SUM[1] ) );
  FA_X1 \intadd_27/U2  ( .A(\intadd_5/SUM[1] ), .B(\intadd_27/B[2] ), .CI(
        \intadd_27/n2 ), .CO(\intadd_27/n1 ), .S(\intadd_16/A[3] ) );
  FA_X1 \intadd_28/U4  ( .A(\intadd_28/A[0] ), .B(\intadd_28/B[0] ), .CI(
        \intadd_28/CI ), .CO(\intadd_28/n3 ), .S(\intadd_28/SUM[0] ) );
  FA_X1 \intadd_28/U3  ( .A(\intadd_28/A[1] ), .B(\intadd_28/B[1] ), .CI(
        \intadd_28/n3 ), .CO(\intadd_28/n2 ), .S(\intadd_28/SUM[1] ) );
  FA_X1 \intadd_28/U2  ( .A(\intadd_28/A[2] ), .B(\intadd_28/B[2] ), .CI(
        \intadd_28/n2 ), .CO(\intadd_28/n1 ), .S(\intadd_28/SUM[2] ) );
  FA_X1 \intadd_29/U4  ( .A(\intadd_29/A[0] ), .B(\intadd_29/B[0] ), .CI(
        \intadd_29/CI ), .CO(\intadd_29/n3 ), .S(\intadd_29/SUM[0] ) );
  FA_X1 \intadd_29/U3  ( .A(\intadd_29/A[1] ), .B(\intadd_29/B[1] ), .CI(
        \intadd_29/n3 ), .CO(\intadd_29/n2 ), .S(\intadd_29/SUM[1] ) );
  FA_X1 \intadd_29/U2  ( .A(\intadd_29/A[2] ), .B(\intadd_19/SUM[0] ), .CI(
        \intadd_29/n2 ), .CO(\intadd_29/n1 ), .S(\intadd_18/B[3] ) );
  FA_X1 \intadd_30/U4  ( .A(\intadd_30/A[0] ), .B(\intadd_30/B[0] ), .CI(
        \intadd_30/CI ), .CO(\intadd_30/n3 ), .S(\intadd_30/SUM[0] ) );
  FA_X1 \intadd_30/U3  ( .A(\intadd_30/A[1] ), .B(\intadd_30/B[1] ), .CI(
        \intadd_30/n3 ), .CO(\intadd_30/n2 ), .S(\intadd_30/SUM[1] ) );
  FA_X1 \intadd_30/U2  ( .A(\intadd_30/A[2] ), .B(\intadd_30/B[2] ), .CI(
        \intadd_30/n2 ), .CO(\intadd_30/n1 ), .S(\intadd_30/SUM[2] ) );
  FA_X1 \intadd_31/U4  ( .A(\intadd_31/A[0] ), .B(\intadd_31/B[0] ), .CI(
        \intadd_9/SUM[0] ), .CO(\intadd_31/n3 ), .S(\intadd_19/A[3] ) );
  FA_X1 \intadd_31/U3  ( .A(\intadd_31/A[1] ), .B(\intadd_9/SUM[1] ), .CI(
        \intadd_31/n3 ), .CO(\intadd_31/n2 ), .S(\intadd_31/SUM[1] ) );
  FA_X1 \intadd_31/U2  ( .A(\intadd_21/SUM[3] ), .B(\intadd_9/SUM[2] ), .CI(
        \intadd_31/n2 ), .CO(\intadd_31/n1 ), .S(\intadd_31/SUM[2] ) );
  FA_X1 \intadd_32/U4  ( .A(\intadd_32/A[0] ), .B(\intadd_32/B[0] ), .CI(
        \intadd_32/CI ), .CO(\intadd_32/n3 ), .S(\intadd_32/SUM[0] ) );
  FA_X1 \intadd_32/U3  ( .A(\intadd_32/A[1] ), .B(\intadd_32/B[1] ), .CI(
        \intadd_32/n3 ), .CO(\intadd_32/n2 ), .S(\intadd_32/SUM[1] ) );
  FA_X1 \intadd_32/U2  ( .A(\intadd_32/A[2] ), .B(\intadd_32/B[2] ), .CI(
        \intadd_32/n2 ), .CO(\intadd_32/n1 ), .S(\intadd_32/SUM[2] ) );
  FA_X1 \intadd_33/U4  ( .A(\intadd_33/A[0] ), .B(\intadd_33/B[0] ), .CI(
        \intadd_33/CI ), .CO(\intadd_33/n3 ), .S(\intadd_33/SUM[0] ) );
  FA_X1 \intadd_33/U3  ( .A(\intadd_7/SUM[0] ), .B(\intadd_33/B[1] ), .CI(
        \intadd_33/n3 ), .CO(\intadd_33/n2 ), .S(\intadd_10/B[3] ) );
  FA_X1 \intadd_33/U2  ( .A(\intadd_33/A[2] ), .B(\intadd_33/B[2] ), .CI(
        \intadd_33/n2 ), .CO(\intadd_33/n1 ), .S(\intadd_10/B[4] ) );
  FA_X1 \intadd_34/U4  ( .A(\intadd_34/A[0] ), .B(\intadd_34/B[0] ), .CI(
        \intadd_34/CI ), .CO(\intadd_34/n3 ), .S(\intadd_32/A[0] ) );
  FA_X1 \intadd_34/U3  ( .A(\intadd_34/A[1] ), .B(\intadd_34/B[1] ), .CI(
        \intadd_34/n3 ), .CO(\intadd_34/n2 ), .S(\intadd_32/B[1] ) );
  FA_X1 \intadd_34/U2  ( .A(\intadd_34/A[2] ), .B(\intadd_34/B[2] ), .CI(
        \intadd_34/n2 ), .CO(\intadd_34/n1 ), .S(\intadd_32/A[2] ) );
  FA_X1 \intadd_35/U4  ( .A(\intadd_35/A[0] ), .B(\intadd_35/B[0] ), .CI(
        \intadd_35/CI ), .CO(\intadd_35/n3 ), .S(\intadd_35/SUM[0] ) );
  FA_X1 \intadd_35/U3  ( .A(\intadd_23/SUM[0] ), .B(\intadd_35/B[1] ), .CI(
        \intadd_35/n3 ), .CO(\intadd_35/n2 ), .S(\intadd_14/B[3] ) );
  FA_X1 \intadd_35/U2  ( .A(\intadd_22/SUM[0] ), .B(\intadd_35/B[2] ), .CI(
        \intadd_35/n2 ), .CO(\intadd_35/n1 ), .S(\intadd_35/SUM[2] ) );
  INV_X1 U1 ( .A(n1201), .ZN(n1132) );
  INV_X1 U2 ( .A(a[1]), .ZN(n1239) );
  NOR2_X2 U3 ( .A1(n565), .A2(n5), .ZN(n1) );
  INV_X2 U4 ( .A(n378), .ZN(n643) );
  NOR2_X1 U5 ( .A1(n1239), .A2(n662), .ZN(n378) );
  NOR2_X2 U8 ( .A1(n726), .A2(n584), .ZN(n717) );
  INV_X1 U9 ( .A(a[15]), .ZN(n84) );
  AND2_X1 U10 ( .A1(n234), .A2(n245), .ZN(n82) );
  OR2_X1 U11 ( .A1(n1238), .A2(n331), .ZN(\intadd_10/A[0] ) );
  INV_X1 U12 ( .A(n337), .ZN(n343) );
  OR2_X1 U13 ( .A1(n950), .A2(n951), .ZN(n974) );
  AND2_X1 U14 ( .A1(n41), .A2(a[11]), .ZN(n817) );
  INV_X1 U15 ( .A(a[9]), .ZN(n767) );
  INV_X1 U16 ( .A(a[11]), .ZN(n480) );
  INV_X1 U17 ( .A(n784), .ZN(n720) );
  INV_X1 U18 ( .A(n817), .ZN(n790) );
  AND2_X1 U19 ( .A1(a[9]), .A2(n179), .ZN(n784) );
  INV_X1 U20 ( .A(a[17]), .ZN(n73) );
  INV_X1 U21 ( .A(n79), .ZN(n776) );
  INV_X1 U22 ( .A(n581), .ZN(n729) );
  AND2_X1 U23 ( .A1(b[0]), .A2(n86), .ZN(n455) );
  INV_X1 U24 ( .A(n54), .ZN(\intadd_29/B[1] ) );
  INV_X1 U25 ( .A(n62), .ZN(\intadd_20/A[1] ) );
  INV_X1 U26 ( .A(n66), .ZN(\intadd_19/A[2] ) );
  INV_X1 U27 ( .A(n106), .ZN(\intadd_10/A[2] ) );
  INV_X1 U28 ( .A(\intadd_32/SUM[0] ), .ZN(\intadd_9/B[3] ) );
  INV_X1 U29 ( .A(n122), .ZN(\intadd_33/A[2] ) );
  AND2_X1 U30 ( .A1(n899), .A2(n900), .ZN(n1017) );
  INV_X1 U31 ( .A(n975), .ZN(n976) );
  OR2_X1 U32 ( .A1(a[7]), .A2(a[8]), .ZN(n356) );
  INV_X1 U33 ( .A(n1147), .ZN(n604) );
  INV_X1 U34 ( .A(n773), .ZN(n774) );
  INV_X1 U35 ( .A(n722), .ZN(n769) );
  AND2_X1 U36 ( .A1(n45), .A2(a[13]), .ZN(\intadd_23/A[0] ) );
  INV_X1 U37 ( .A(n82), .ZN(n690) );
  INV_X1 U38 ( .A(n71), .ZN(n77) );
  INV_X1 U39 ( .A(n36), .ZN(n37) );
  INV_X1 U40 ( .A(n449), .ZN(n38) );
  INV_X1 U41 ( .A(n317), .ZN(n410) );
  AND2_X1 U42 ( .A1(a[13]), .A2(n52), .ZN(n246) );
  AND2_X1 U43 ( .A1(a[17]), .A2(n86), .ZN(n845) );
  INV_X1 U44 ( .A(a[20]), .ZN(n156) );
  INV_X1 U45 ( .A(a[19]), .ZN(n842) );
  INV_X1 U46 ( .A(a[7]), .ZN(n772) );
  AND2_X1 U47 ( .A1(n260), .A2(a[11]), .ZN(n818) );
  AND2_X1 U48 ( .A1(b[0]), .A2(n52), .ZN(n495) );
  INV_X1 U49 ( .A(n447), .ZN(n448) );
  INV_X1 U50 ( .A(n88), .ZN(\intadd_21/A[1] ) );
  INV_X1 U51 ( .A(n100), .ZN(\intadd_10/A[1] ) );
  INV_X1 U52 ( .A(n409), .ZN(n318) );
  INV_X1 U53 ( .A(n338), .ZN(n339) );
  OR2_X1 U54 ( .A1(\intadd_5/SUM[2] ), .A2(n937), .ZN(n938) );
  AND2_X1 U55 ( .A1(n829), .A2(a[9]), .ZN(n830) );
  OR2_X1 U56 ( .A1(n268), .A2(n267), .ZN(n281) );
  INV_X1 U57 ( .A(\intadd_4/SUM[4] ), .ZN(n950) );
  INV_X1 U58 ( .A(n845), .ZN(n825) );
  AND2_X1 U59 ( .A1(n74), .A2(a[17]), .ZN(n984) );
  INV_X1 U60 ( .A(n1096), .ZN(n1104) );
  INV_X1 U61 ( .A(n626), .ZN(n1103) );
  INV_X1 U62 ( .A(n1150), .ZN(n1138) );
  INV_X1 U63 ( .A(a[21]), .ZN(n1095) );
  INV_X1 U64 ( .A(n624), .ZN(n1101) );
  INV_X1 U65 ( .A(n373), .ZN(n661) );
  INV_X1 U66 ( .A(a[3]), .ZN(n565) );
  INV_X1 U67 ( .A(n21), .ZN(n93) );
  INV_X1 U68 ( .A(n18), .ZN(n519) );
  INV_X1 U69 ( .A(n192), .ZN(n201) );
  INV_X1 U70 ( .A(n58), .ZN(\intadd_29/A[2] ) );
  OR2_X1 U71 ( .A1(n1000), .A2(n397), .ZN(n925) );
  INV_X1 U72 ( .A(\intadd_34/n1 ), .ZN(\intadd_7/A[2] ) );
  AND2_X1 U73 ( .A1(n102), .A2(a[19]), .ZN(\intadd_12/A[1] ) );
  INV_X1 U74 ( .A(n1141), .ZN(n1108) );
  INV_X1 U75 ( .A(b[23]), .ZN(n1151) );
  INV_X1 U76 ( .A(b[0]), .ZN(n1238) );
  AND2_X1 U77 ( .A1(n522), .A2(n521), .ZN(n537) );
  INV_X1 U78 ( .A(n193), .ZN(n1053) );
  INV_X1 U79 ( .A(n1050), .ZN(n1054) );
  INV_X1 U80 ( .A(n205), .ZN(n206) );
  INV_X1 U81 ( .A(n29), .ZN(\intadd_8/A[1] ) );
  INV_X1 U82 ( .A(\intadd_0/SUM[1] ), .ZN(n542) );
  INV_X1 U83 ( .A(n182), .ZN(n183) );
  INV_X1 U84 ( .A(\intadd_30/SUM[0] ), .ZN(\intadd_20/A[3] ) );
  INV_X1 U85 ( .A(\intadd_30/SUM[2] ), .ZN(n1212) );
  INV_X1 U86 ( .A(\intadd_30/SUM[1] ), .ZN(\intadd_19/B[3] ) );
  INV_X1 U87 ( .A(\intadd_32/SUM[1] ), .ZN(\intadd_9/B[4] ) );
  INV_X1 U88 ( .A(\intadd_32/SUM[2] ), .ZN(\intadd_10/A[4] ) );
  INV_X1 U89 ( .A(n1002), .ZN(n1073) );
  INV_X1 U90 ( .A(n934), .ZN(n940) );
  INV_X1 U91 ( .A(n997), .ZN(n1084) );
  INV_X1 U92 ( .A(n1177), .ZN(n960) );
  INV_X1 U93 ( .A(n1255), .ZN(n1023) );
  INV_X1 U94 ( .A(n1202), .ZN(n1065) );
  INV_X1 U95 ( .A(n153), .ZN(\intadd_2/B[4] ) );
  INV_X1 U96 ( .A(n1164), .ZN(n1162) );
  INV_X1 U97 ( .A(b[23]), .ZN(n1163) );
  INV_X1 U98 ( .A(a[0]), .ZN(n1246) );
  INV_X1 U99 ( .A(b[0]), .ZN(n1247) );
  INV_X1 U100 ( .A(n1279), .ZN(n1276) );
  INV_X1 U101 ( .A(\intadd_28/n1 ), .ZN(\intadd_0/B[4] ) );
  INV_X1 U102 ( .A(n995), .ZN(n1194) );
  INV_X1 U103 ( .A(n1268), .ZN(n1270) );
  INV_X1 U104 ( .A(n1264), .ZN(n1266) );
  INV_X1 U105 ( .A(n1226), .ZN(n1014) );
  NOR2_X2 U106 ( .A1(a[3]), .A2(n5), .ZN(n633) );
  INV_X1 U107 ( .A(b[16]), .ZN(n575) );
  INV_X1 U108 ( .A(b[22]), .ZN(n1140) );
  INV_X1 U109 ( .A(b[12]), .ZN(n650) );
  INV_X1 U110 ( .A(b[18]), .ZN(n1114) );
  INV_X1 U111 ( .A(b[2]), .ZN(n606) );
  INV_X1 U112 ( .A(b[8]), .ZN(n654) );
  INV_X1 U113 ( .A(b[15]), .ZN(n687) );
  INV_X1 U114 ( .A(b[21]), .ZN(n878) );
  INV_X1 U115 ( .A(b[19]), .ZN(n1106) );
  INV_X1 U116 ( .A(b[7]), .ZN(n712) );
  INV_X1 U117 ( .A(b[9]), .ZN(n689) );
  INV_X1 U118 ( .A(n305), .ZN(n92) );
  INV_X1 U119 ( .A(n569), .ZN(n570) );
  INV_X1 U120 ( .A(n735), .ZN(n740) );
  INV_X1 U121 ( .A(n174), .ZN(n168) );
  INV_X1 U122 ( .A(n315), .ZN(n417) );
  INV_X1 U123 ( .A(n636), .ZN(n367) );
  INV_X1 U124 ( .A(n585), .ZN(n663) );
  INV_X1 U125 ( .A(n768), .ZN(n179) );
  INV_X1 U126 ( .A(n145), .ZN(n147) );
  INV_X1 U127 ( .A(n747), .ZN(n144) );
  INV_X1 U128 ( .A(n691), .ZN(n235) );
  INV_X1 U129 ( .A(a[6]), .ZN(n20) );
  INV_X1 U130 ( .A(n530), .ZN(n508) );
  INV_X1 U131 ( .A(a[13]), .ZN(n245) );
  INV_X1 U132 ( .A(b[11]), .ZN(n754) );
  INV_X1 U133 ( .A(n246), .ZN(n812) );
  INV_X1 U134 ( .A(b[13]), .ZN(n637) );
  INV_X1 U135 ( .A(\intadd_9/SUM[4] ), .ZN(n904) );
  INV_X1 U136 ( .A(n576), .ZN(n701) );
  INV_X1 U137 ( .A(n605), .ZN(n369) );
  INV_X1 U138 ( .A(n668), .ZN(n666) );
  INV_X1 U139 ( .A(n514), .ZN(n584) );
  INV_X1 U140 ( .A(n795), .ZN(n148) );
  INV_X1 U141 ( .A(b[14]), .ZN(n554) );
  INV_X1 U142 ( .A(b[17]), .ZN(n824) );
  INV_X1 U143 ( .A(n207), .ZN(n204) );
  INV_X1 U144 ( .A(b[5]), .ZN(n741) );
  INV_X1 U145 ( .A(b[1]), .ZN(n628) );
  INV_X1 U146 ( .A(b[6]), .ZN(n764) );
  INV_X1 U147 ( .A(b[4]), .ZN(n704) );
  INV_X1 U148 ( .A(n469), .ZN(n471) );
  INV_X1 U149 ( .A(n400), .ZN(n320) );
  INV_X1 U150 ( .A(n385), .ZN(n345) );
  INV_X1 U151 ( .A(n384), .ZN(n386) );
  INV_X1 U152 ( .A(n970), .ZN(n966) );
  INV_X1 U153 ( .A(n623), .ZN(n1100) );
  INV_X1 U154 ( .A(b[3]), .ZN(n555) );
  INV_X1 U155 ( .A(b[10]), .ZN(n649) );
  INV_X1 U156 ( .A(n472), .ZN(n450) );
  INV_X1 U157 ( .A(n902), .ZN(n903) );
  INV_X1 U158 ( .A(\intadd_5/SUM[3] ), .ZN(n944) );
  INV_X1 U159 ( .A(n1181), .ZN(n972) );
  INV_X1 U160 ( .A(n1133), .ZN(n973) );
  INV_X1 U161 ( .A(b[20]), .ZN(n1098) );
  INV_X1 U162 ( .A(n1092), .ZN(n1007) );
  INV_X1 U163 ( .A(n1020), .ZN(n1021) );
  INV_X1 U164 ( .A(n1028), .ZN(n1034) );
  INV_X1 U165 ( .A(n1047), .ZN(n1045) );
  INV_X1 U166 ( .A(n1089), .ZN(n1091) );
  INV_X1 U167 ( .A(n1010), .ZN(n1256) );
  INV_X1 U168 ( .A(n1061), .ZN(n1063) );
  INV_X1 U169 ( .A(n1033), .ZN(n1029) );
  INV_X1 U170 ( .A(n1248), .ZN(n1035) );
  INV_X1 U171 ( .A(n1225), .ZN(n981) );
  INV_X1 U172 ( .A(n1230), .ZN(n1232) );
  INV_X1 U173 ( .A(n1231), .ZN(n1137) );
  INV_X1 U174 ( .A(n1195), .ZN(n1179) );
  NAND2_X1 U175 ( .A1(a[0]), .A2(a[1]), .ZN(n527) );
  NAND2_X1 U176 ( .A1(a[0]), .A2(n1239), .ZN(n528) );
  NOR2_X1 U177 ( .A1(a[0]), .A2(n1239), .ZN(n530) );
  NAND2_X1 U178 ( .A1(n530), .A2(n628), .ZN(n2) );
  OAI221_X1 U179 ( .B1(b[2]), .B2(n527), .C1(n606), .C2(n528), .A(n2), .ZN(
        n1041) );
  NOR2_X1 U180 ( .A1(a[1]), .A2(a[2]), .ZN(n373) );
  NAND2_X1 U181 ( .A1(a[1]), .A2(a[2]), .ZN(n376) );
  NAND2_X1 U182 ( .A1(n661), .A2(n376), .ZN(n5) );
  OAI21_X1 U183 ( .B1(n628), .B2(n1246), .A(a[1]), .ZN(n3) );
  AOI22_X1 U184 ( .A1(b[0]), .A2(n5), .B1(n3), .B2(n1247), .ZN(n1040) );
  NAND2_X1 U185 ( .A1(n1041), .A2(n1040), .ZN(n1275) );
  OAI211_X1 U186 ( .C1(n373), .C2(n1238), .A(n376), .B(a[3]), .ZN(n1274) );
  NAND2_X1 U187 ( .A1(n530), .A2(n606), .ZN(n4) );
  OAI221_X1 U188 ( .B1(b[3]), .B2(n527), .C1(n555), .C2(n528), .A(n4), .ZN(n8)
         );
  NAND2_X1 U189 ( .A1(a[3]), .A2(n373), .ZN(n631) );
  NAND2_X1 U190 ( .A1(n565), .A2(a[2]), .ZN(n662) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(n633), .B1(n1), .B2(n628), .ZN(n6) );
  OAI221_X1 U192 ( .B1(b[0]), .B2(n631), .C1(n1238), .C2(n643), .A(n6), .ZN(n7) );
  NAND2_X1 U193 ( .A1(n8), .A2(n7), .ZN(n1277) );
  INV_X1 U194 ( .A(n1277), .ZN(n1278) );
  NOR2_X1 U195 ( .A1(n8), .A2(n7), .ZN(n534) );
  OR2_X1 U196 ( .A1(n1278), .A2(n534), .ZN(n1273) );
  FA_X1 U197 ( .A(\intadd_20/SUM[2] ), .B(\intadd_19/SUM[1] ), .CI(
        \intadd_29/n1 ), .CO(n1216), .S(n1219) );
  AOI22_X1 U198 ( .A1(n1216), .A2(\intadd_20/SUM[3] ), .B1(n1219), .B2(
        \intadd_18/n1 ), .ZN(n910) );
  INV_X2 U199 ( .A(\intadd_0/n1 ), .ZN(n909) );
  AND3_X1 U200 ( .A1(\intadd_20/SUM[2] ), .A2(\intadd_29/n1 ), .A3(
        \intadd_19/SUM[1] ), .ZN(n10) );
  NOR3_X1 U201 ( .A1(\intadd_20/SUM[3] ), .A2(\intadd_18/n1 ), .A3(n10), .ZN(
        n908) );
  NOR4_X1 U202 ( .A1(\intadd_18/n1 ), .A2(\intadd_20/SUM[2] ), .A3(
        \intadd_29/n1 ), .A4(\intadd_19/SUM[1] ), .ZN(n11) );
  NOR2_X1 U203 ( .A1(n1216), .A2(\intadd_20/SUM[3] ), .ZN(n1215) );
  NOR2_X1 U204 ( .A1(n11), .A2(n1215), .ZN(n912) );
  INV_X1 U205 ( .A(n912), .ZN(n12) );
  AOI211_X1 U206 ( .C1(n910), .C2(n909), .A(n908), .B(n12), .ZN(n1207) );
  INV_X2 U207 ( .A(n13), .ZN(\d[18] ) );
  INV_X2 U208 ( .A(\intadd_11/SUM[0] ), .ZN(\d[20] ) );
  INV_X2 U209 ( .A(\intadd_11/SUM[1] ), .ZN(\d[21] ) );
  INV_X2 U210 ( .A(\intadd_8/n1 ), .ZN(\intadd_0/B[3] ) );
  AND2_X2 U211 ( .A1(a[3]), .A2(a[4]), .ZN(n580) );
  INV_X2 U212 ( .A(a[5]), .ZN(n726) );
  NOR2_X1 U213 ( .A1(n580), .A2(n726), .ZN(\intadd_3/B[0] ) );
  AOI221_X1 U214 ( .B1(a[1]), .B2(b[7]), .C1(n1239), .C2(n712), .A(n1246), 
        .ZN(n14) );
  AOI21_X1 U215 ( .B1(n530), .B2(n764), .A(n14), .ZN(n188) );
  NAND2_X1 U216 ( .A1(n726), .A2(n580), .ZN(n581) );
  NOR2_X1 U217 ( .A1(a[3]), .A2(a[4]), .ZN(n514) );
  NOR2_X1 U218 ( .A1(n580), .A2(n514), .ZN(n526) );
  NAND2_X1 U219 ( .A1(n526), .A2(n726), .ZN(n715) );
  AND2_X2 U220 ( .A1(\intadd_3/B[0] ), .A2(n584), .ZN(n727) );
  INV_X2 U221 ( .A(n727), .ZN(n714) );
  AOI22_X1 U222 ( .A1(b[3]), .A2(n715), .B1(n714), .B2(n555), .ZN(n15) );
  AOI221_X1 U223 ( .B1(n729), .B2(b[2]), .C1(n717), .C2(n606), .A(n15), .ZN(
        n187) );
  AOI22_X1 U224 ( .A1(b[4]), .A2(n643), .B1(n631), .B2(n704), .ZN(n16) );
  AOI221_X1 U225 ( .B1(n633), .B2(b[5]), .C1(n1), .C2(n741), .A(n16), .ZN(n186) );
  AOI22_X1 U226 ( .A1(a[5]), .A2(a[6]), .B1(n20), .B2(n726), .ZN(n21) );
  NOR2_X1 U227 ( .A1(n93), .A2(n1238), .ZN(n540) );
  AOI22_X1 U228 ( .A1(b[6]), .A2(n528), .B1(n527), .B2(n764), .ZN(n17) );
  AOI21_X1 U229 ( .B1(n530), .B2(n741), .A(n17), .ZN(n18) );
  AOI22_X1 U230 ( .A1(b[1]), .A2(n729), .B1(n717), .B2(n628), .ZN(n19) );
  OAI221_X1 U231 ( .B1(b[2]), .B2(n714), .C1(n606), .C2(n715), .A(n19), .ZN(
        n518) );
  AOI222_X1 U232 ( .A1(n540), .A2(n519), .B1(n540), .B2(n518), .C1(n519), .C2(
        n518), .ZN(n196) );
  NOR2_X1 U233 ( .A1(n726), .A2(n20), .ZN(n22) );
  NOR2_X1 U234 ( .A1(n22), .A2(n772), .ZN(n761) );
  NOR3_X1 U235 ( .A1(a[5]), .A2(a[6]), .A3(n772), .ZN(n725) );
  AOI21_X1 U236 ( .B1(n761), .B2(n628), .A(n725), .ZN(n505) );
  NAND2_X1 U237 ( .A1(a[7]), .A2(n21), .ZN(n773) );
  NAND2_X1 U238 ( .A1(n21), .A2(n772), .ZN(n723) );
  OAI22_X1 U239 ( .A1(b[0]), .A2(n773), .B1(n723), .B2(n628), .ZN(n24) );
  NAND2_X1 U240 ( .A1(n772), .A2(n22), .ZN(n79) );
  AOI21_X1 U241 ( .B1(n79), .B2(n505), .A(n1247), .ZN(n23) );
  AOI21_X1 U242 ( .B1(n505), .B2(n24), .A(n23), .ZN(n195) );
  INV_X2 U243 ( .A(n25), .ZN(\intadd_26/A[2] ) );
  AOI22_X1 U244 ( .A1(b[3]), .A2(n723), .B1(n773), .B2(n555), .ZN(n26) );
  AOI221_X1 U245 ( .B1(n776), .B2(b[2]), .C1(n725), .C2(n606), .A(n26), .ZN(
        n166) );
  AOI22_X1 U246 ( .A1(b[5]), .A2(n715), .B1(n714), .B2(n741), .ZN(n27) );
  AOI221_X1 U247 ( .B1(n729), .B2(b[4]), .C1(n717), .C2(n704), .A(n27), .ZN(
        n165) );
  AOI22_X1 U248 ( .A1(b[6]), .A2(n643), .B1(n631), .B2(n764), .ZN(n28) );
  AOI221_X1 U249 ( .B1(n633), .B2(b[7]), .C1(n1), .C2(n712), .A(n28), .ZN(n164) );
  INV_X2 U250 ( .A(\intadd_0/SUM[2] ), .ZN(\intadd_8/A[4] ) );
  NOR2_X1 U251 ( .A1(a[9]), .A2(a[10]), .ZN(n497) );
  AOI21_X1 U252 ( .B1(a[10]), .B2(a[9]), .A(n497), .ZN(n41) );
  NAND2_X1 U253 ( .A1(b[0]), .A2(n41), .ZN(n167) );
  NAND2_X1 U254 ( .A1(a[7]), .A2(a[8]), .ZN(n829) );
  NOR2_X1 U255 ( .A1(a[9]), .A2(n829), .ZN(n771) );
  NOR3_X1 U256 ( .A1(a[7]), .A2(a[8]), .A3(n767), .ZN(n722) );
  NAND2_X1 U257 ( .A1(n829), .A2(n356), .ZN(n768) );
  NAND2_X1 U258 ( .A1(n179), .A2(n767), .ZN(n780) );
  AOI22_X1 U259 ( .A1(b[2]), .A2(n780), .B1(n720), .B2(n606), .ZN(n30) );
  AOI221_X1 U260 ( .B1(n771), .B2(b[1]), .C1(n722), .C2(n628), .A(n30), .ZN(
        n170) );
  AOI22_X1 U261 ( .A1(b[4]), .A2(n723), .B1(n773), .B2(n704), .ZN(n31) );
  AOI221_X1 U262 ( .B1(n776), .B2(b[3]), .C1(n725), .C2(n555), .A(n31), .ZN(
        n173) );
  OAI21_X1 U263 ( .B1(n170), .B2(n167), .A(n173), .ZN(n32) );
  INV_X2 U264 ( .A(n32), .ZN(n33) );
  AOI21_X1 U265 ( .B1(n167), .B2(n170), .A(n33), .ZN(n34) );
  INV_X2 U266 ( .A(n34), .ZN(\intadd_0/A[1] ) );
  INV_X2 U267 ( .A(\intadd_28/SUM[1] ), .ZN(\intadd_0/A[2] ) );
  INV_X2 U268 ( .A(\intadd_28/SUM[2] ), .ZN(\intadd_0/A[3] ) );
  INV_X2 U269 ( .A(\intadd_29/SUM[0] ), .ZN(\intadd_28/B[1] ) );
  INV_X2 U270 ( .A(\intadd_18/SUM[2] ), .ZN(\intadd_28/B[2] ) );
  INV_X2 U271 ( .A(\intadd_29/SUM[1] ), .ZN(\intadd_28/A[2] ) );
  NAND2_X1 U272 ( .A1(a[13]), .A2(a[14]), .ZN(n35) );
  OAI21_X1 U273 ( .B1(a[13]), .B2(a[14]), .A(n35), .ZN(n83) );
  NOR2_X1 U274 ( .A1(a[15]), .A2(n83), .ZN(n694) );
  NOR2_X1 U275 ( .A1(a[14]), .A2(n84), .ZN(n234) );
  AOI21_X1 U276 ( .B1(a[13]), .B2(a[14]), .A(n84), .ZN(n288) );
  OAI21_X1 U277 ( .B1(n1247), .B2(n628), .A(n288), .ZN(n36) );
  AOI211_X1 U278 ( .C1(b[1]), .C2(n694), .A(n82), .B(n37), .ZN(n39) );
  NAND3_X1 U279 ( .A1(a[13]), .A2(a[14]), .A3(n84), .ZN(n691) );
  OAI211_X1 U280 ( .C1(n628), .C2(n82), .A(n1247), .B(n288), .ZN(n449) );
  AOI221_X1 U281 ( .B1(n1238), .B2(n39), .C1(n691), .C2(n39), .A(n38), .ZN(n65) );
  NOR2_X1 U282 ( .A1(a[12]), .A2(a[11]), .ZN(n47) );
  AOI21_X1 U283 ( .B1(a[11]), .B2(a[12]), .A(n47), .ZN(n52) );
  NAND2_X1 U284 ( .A1(n52), .A2(n245), .ZN(n813) );
  NAND2_X1 U285 ( .A1(a[12]), .A2(a[11]), .ZN(n45) );
  NOR2_X1 U286 ( .A1(a[13]), .A2(n45), .ZN(n816) );
  NOR3_X1 U287 ( .A1(a[12]), .A2(a[11]), .A3(n245), .ZN(n815) );
  AOI22_X1 U288 ( .A1(b[1]), .A2(n816), .B1(n815), .B2(n628), .ZN(n40) );
  OAI221_X1 U289 ( .B1(b[2]), .B2(n812), .C1(n606), .C2(n813), .A(n40), .ZN(
        n61) );
  NOR2_X1 U290 ( .A1(n1247), .A2(n83), .ZN(n60) );
  NAND2_X1 U291 ( .A1(n41), .A2(n480), .ZN(n791) );
  NAND2_X1 U292 ( .A1(a[9]), .A2(a[10]), .ZN(n260) );
  NOR2_X1 U293 ( .A1(a[11]), .A2(n260), .ZN(n819) );
  AOI22_X1 U294 ( .A1(b[3]), .A2(n819), .B1(n793), .B2(n555), .ZN(n42) );
  OAI221_X1 U295 ( .B1(b[4]), .B2(n790), .C1(n704), .C2(n791), .A(n42), .ZN(
        n59) );
  AOI22_X1 U296 ( .A1(b[13]), .A2(n633), .B1(n1), .B2(n637), .ZN(n43) );
  OAI221_X1 U297 ( .B1(b[12]), .B2(n631), .C1(n650), .C2(n643), .A(n43), .ZN(
        n63) );
  INV_X2 U298 ( .A(n44), .ZN(\intadd_20/B[2] ) );
  AOI22_X1 U299 ( .A1(b[1]), .A2(n813), .B1(n812), .B2(n628), .ZN(n46) );
  AOI221_X1 U300 ( .B1(n816), .B2(b[0]), .C1(n815), .C2(n1238), .A(n46), .ZN(
        n490) );
  OAI21_X1 U301 ( .B1(n47), .B2(n1247), .A(\intadd_23/A[0] ), .ZN(n489) );
  NOR2_X1 U302 ( .A1(n490), .A2(n489), .ZN(n57) );
  AOI22_X1 U303 ( .A1(b[9]), .A2(n729), .B1(n717), .B2(n689), .ZN(n48) );
  OAI221_X1 U304 ( .B1(b[10]), .B2(n714), .C1(n649), .C2(n715), .A(n48), .ZN(
        n56) );
  AOI22_X1 U305 ( .A1(b[12]), .A2(n633), .B1(n1), .B2(n650), .ZN(n49) );
  OAI221_X1 U306 ( .B1(b[11]), .B2(n631), .C1(n754), .C2(n643), .A(n49), .ZN(
        n55) );
  INV_X2 U307 ( .A(n50), .ZN(\intadd_20/A[2] ) );
  AOI22_X1 U308 ( .A1(b[3]), .A2(n771), .B1(n722), .B2(n555), .ZN(n51) );
  OAI221_X1 U309 ( .B1(b[4]), .B2(n720), .C1(n704), .C2(n780), .A(n51), .ZN(
        n496) );
  AOI22_X1 U310 ( .A1(b[1]), .A2(n819), .B1(n793), .B2(n628), .ZN(n53) );
  OAI221_X1 U311 ( .B1(b[2]), .B2(n790), .C1(n606), .C2(n791), .A(n53), .ZN(
        n494) );
  FA_X1 U312 ( .A(n57), .B(n56), .CI(n55), .CO(n50), .S(n58) );
  FA_X1 U313 ( .A(n61), .B(n60), .CI(n59), .CO(n64), .S(n62) );
  FA_X1 U314 ( .A(n65), .B(n64), .CI(n63), .CO(n66), .S(n44) );
  INV_X2 U315 ( .A(\intadd_21/SUM[0] ), .ZN(\intadd_30/CI ) );
  AOI22_X1 U316 ( .A1(b[8]), .A2(n780), .B1(n720), .B2(n654), .ZN(n67) );
  AOI221_X1 U317 ( .B1(n771), .B2(b[7]), .C1(n722), .C2(n712), .A(n67), .ZN(
        n453) );
  AOI22_X1 U318 ( .A1(b[6]), .A2(n791), .B1(n790), .B2(n764), .ZN(n68) );
  AOI221_X1 U319 ( .B1(n819), .B2(b[5]), .C1(n793), .C2(n741), .A(n68), .ZN(
        n452) );
  AOI221_X1 U320 ( .B1(b[16]), .B2(a[1]), .C1(n575), .C2(n1239), .A(n1246), 
        .ZN(n69) );
  AOI21_X1 U321 ( .B1(n530), .B2(n687), .A(n69), .ZN(n451) );
  INV_X2 U322 ( .A(n70), .ZN(\intadd_30/A[0] ) );
  NOR3_X1 U323 ( .A1(a[15]), .A2(a[16]), .A3(n73), .ZN(n828) );
  NAND2_X1 U324 ( .A1(a[15]), .A2(a[16]), .ZN(n74) );
  OAI21_X1 U325 ( .B1(n1247), .B2(n828), .A(n984), .ZN(n71) );
  NOR2_X1 U326 ( .A1(a[15]), .A2(a[16]), .ZN(n72) );
  AOI21_X1 U327 ( .B1(a[16]), .B2(a[15]), .A(n72), .ZN(n86) );
  NAND2_X1 U328 ( .A1(n86), .A2(n73), .ZN(n826) );
  NOR2_X1 U329 ( .A1(a[17]), .A2(n74), .ZN(n846) );
  AOI21_X1 U330 ( .B1(n846), .B2(b[0]), .A(n828), .ZN(n75) );
  OAI221_X1 U331 ( .B1(b[1]), .B2(n825), .C1(n628), .C2(n826), .A(n75), .ZN(
        n76) );
  NAND3_X1 U332 ( .A1(n1238), .A2(n76), .A3(n984), .ZN(n436) );
  OAI21_X1 U333 ( .B1(n77), .B2(n76), .A(n436), .ZN(n459) );
  AOI22_X1 U334 ( .A1(b[13]), .A2(n715), .B1(n714), .B2(n637), .ZN(n78) );
  AOI221_X1 U335 ( .B1(n729), .B2(b[12]), .C1(n717), .C2(n650), .A(n78), .ZN(
        n458) );
  AOI22_X1 U336 ( .A1(a[7]), .A2(n754), .B1(b[11]), .B2(n772), .ZN(n94) );
  OAI22_X1 U337 ( .A1(n79), .A2(n649), .B1(n93), .B2(n94), .ZN(n80) );
  AOI21_X1 U338 ( .B1(n725), .B2(n649), .A(n80), .ZN(n457) );
  INV_X2 U339 ( .A(n81), .ZN(\intadd_30/B[1] ) );
  INV_X2 U340 ( .A(\intadd_21/SUM[1] ), .ZN(\intadd_30/A[1] ) );
  INV_X2 U341 ( .A(\intadd_31/SUM[1] ), .ZN(\intadd_30/B[2] ) );
  INV_X2 U342 ( .A(\intadd_21/SUM[2] ), .ZN(\intadd_30/A[2] ) );
  NOR2_X1 U343 ( .A1(n84), .A2(n83), .ZN(n693) );
  AOI22_X1 U344 ( .A1(b[2]), .A2(n694), .B1(n693), .B2(n606), .ZN(n85) );
  OAI221_X1 U345 ( .B1(b[1]), .B2(n690), .C1(n628), .C2(n691), .A(n85), .ZN(
        n456) );
  AOI22_X1 U346 ( .A1(b[3]), .A2(n816), .B1(n815), .B2(n555), .ZN(n87) );
  OAI221_X1 U347 ( .B1(b[4]), .B2(n812), .C1(n704), .C2(n813), .A(n87), .ZN(
        n454) );
  AOI22_X1 U348 ( .A1(b[16]), .A2(n633), .B1(n1), .B2(n575), .ZN(n89) );
  OAI221_X1 U349 ( .B1(b[15]), .B2(n631), .C1(n687), .C2(n643), .A(n89), .ZN(
        n99) );
  AOI22_X1 U350 ( .A1(a[9]), .A2(n689), .B1(b[9]), .B2(n767), .ZN(n429) );
  AOI221_X1 U351 ( .B1(a[8]), .B2(n689), .C1(n772), .C2(b[9]), .A(n429), .ZN(
        n90) );
  OAI22_X1 U352 ( .A1(n179), .A2(n90), .B1(b[10]), .B2(n780), .ZN(n91) );
  AOI21_X1 U353 ( .B1(n784), .B2(b[10]), .A(n91), .ZN(n98) );
  NOR2_X1 U354 ( .A1(n776), .A2(n725), .ZN(n95) );
  AOI22_X1 U355 ( .A1(a[7]), .A2(b[12]), .B1(n650), .B2(n772), .ZN(n305) );
  OAI22_X1 U356 ( .A1(n95), .A2(n94), .B1(n93), .B2(n92), .ZN(n97) );
  INV_X2 U357 ( .A(n96), .ZN(\intadd_9/B[1] ) );
  FA_X1 U358 ( .A(n99), .B(n98), .CI(n97), .CO(n100), .S(n96) );
  NAND2_X1 U359 ( .A1(a[17]), .A2(a[18]), .ZN(n102) );
  AOI22_X1 U360 ( .A1(b[15]), .A2(n729), .B1(n717), .B2(n687), .ZN(n101) );
  OAI221_X1 U361 ( .B1(b[16]), .B2(n714), .C1(n575), .C2(n715), .A(n101), .ZN(
        n113) );
  OAI21_X1 U362 ( .B1(a[17]), .B2(a[18]), .A(n102), .ZN(n331) );
  NOR2_X1 U363 ( .A1(a[19]), .A2(n331), .ZN(n882) );
  NOR2_X1 U364 ( .A1(n842), .A2(n331), .ZN(n881) );
  NAND3_X1 U365 ( .A1(a[17]), .A2(a[18]), .A3(n842), .ZN(n884) );
  NOR2_X1 U366 ( .A1(a[17]), .A2(a[18]), .ZN(n104) );
  NAND2_X1 U367 ( .A1(a[19]), .A2(n104), .ZN(n885) );
  AOI22_X1 U368 ( .A1(b[0]), .A2(n884), .B1(n885), .B2(n1247), .ZN(n103) );
  AOI221_X1 U369 ( .B1(n882), .B2(b[1]), .C1(n881), .C2(n628), .A(n103), .ZN(
        n330) );
  OAI21_X1 U370 ( .B1(n104), .B2(n1247), .A(\intadd_12/A[1] ), .ZN(n329) );
  NOR2_X1 U371 ( .A1(n330), .A2(n329), .ZN(n112) );
  AOI22_X1 U372 ( .A1(b[13]), .A2(n776), .B1(n725), .B2(n637), .ZN(n105) );
  OAI221_X1 U373 ( .B1(b[14]), .B2(n773), .C1(n554), .C2(n723), .A(n105), .ZN(
        n111) );
  AOI22_X1 U374 ( .A1(b[15]), .A2(n723), .B1(n773), .B2(n687), .ZN(n107) );
  AOI221_X1 U375 ( .B1(n776), .B2(b[14]), .C1(n725), .C2(n554), .A(n107), .ZN(
        n342) );
  AOI22_X1 U376 ( .A1(b[6]), .A2(n691), .B1(n690), .B2(n764), .ZN(n108) );
  AOI221_X1 U377 ( .B1(n694), .B2(b[7]), .C1(n693), .C2(n712), .A(n108), .ZN(
        n341) );
  AOI22_X1 U378 ( .A1(b[17]), .A2(n715), .B1(n714), .B2(n824), .ZN(n109) );
  AOI221_X1 U379 ( .B1(n729), .B2(b[16]), .C1(n717), .C2(n575), .A(n109), .ZN(
        n340) );
  INV_X2 U380 ( .A(n110), .ZN(n121) );
  FA_X1 U381 ( .A(n113), .B(n112), .CI(n111), .CO(n120), .S(n106) );
  AOI22_X1 U382 ( .A1(b[11]), .A2(n791), .B1(n790), .B2(n754), .ZN(n114) );
  AOI221_X1 U383 ( .B1(n819), .B2(b[10]), .C1(n793), .C2(n649), .A(n114), .ZN(
        n348) );
  AOI22_X1 U384 ( .A1(b[21]), .A2(n528), .B1(n527), .B2(n878), .ZN(n115) );
  AOI21_X1 U385 ( .B1(n530), .B2(n1098), .A(n115), .ZN(n347) );
  AOI22_X1 U386 ( .A1(b[18]), .A2(n643), .B1(n631), .B2(n1114), .ZN(n116) );
  AOI221_X1 U387 ( .B1(n633), .B2(b[19]), .C1(n1), .C2(n1106), .A(n116), .ZN(
        n346) );
  INV_X2 U388 ( .A(n117), .ZN(n119) );
  INV_X2 U389 ( .A(n118), .ZN(\intadd_10/A[3] ) );
  FA_X1 U390 ( .A(n121), .B(n120), .CI(n119), .CO(n122), .S(n118) );
  AOI22_X1 U391 ( .A1(b[20]), .A2(n528), .B1(n527), .B2(n1098), .ZN(n123) );
  AOI21_X1 U392 ( .B1(n530), .B2(n1106), .A(n123), .ZN(n336) );
  AOI22_X1 U393 ( .A1(b[8]), .A2(n813), .B1(n812), .B2(n654), .ZN(n124) );
  AOI221_X1 U394 ( .B1(n816), .B2(b[7]), .C1(n815), .C2(n712), .A(n124), .ZN(
        n335) );
  AOI22_X1 U395 ( .A1(b[5]), .A2(n691), .B1(n690), .B2(n741), .ZN(n125) );
  AOI221_X1 U396 ( .B1(n694), .B2(b[6]), .C1(n693), .C2(n764), .A(n125), .ZN(
        n334) );
  INV_X2 U397 ( .A(n126), .ZN(\intadd_32/CI ) );
  INV_X2 U398 ( .A(\intadd_33/SUM[0] ), .ZN(\intadd_32/B[0] ) );
  INV_X2 U399 ( .A(\intadd_7/SUM[1] ), .ZN(\intadd_32/B[2] ) );
  AOI22_X1 U400 ( .A1(b[10]), .A2(n813), .B1(n812), .B2(n649), .ZN(n127) );
  AOI221_X1 U401 ( .B1(n816), .B2(b[9]), .C1(n815), .C2(n689), .A(n127), .ZN(
        n352) );
  AOI22_X1 U402 ( .A1(b[12]), .A2(n791), .B1(n790), .B2(n650), .ZN(n128) );
  AOI221_X1 U403 ( .B1(n819), .B2(b[11]), .C1(n793), .C2(n754), .A(n128), .ZN(
        n351) );
  AOI22_X1 U404 ( .A1(b[19]), .A2(n643), .B1(n631), .B2(n1106), .ZN(n129) );
  AOI221_X1 U405 ( .B1(n633), .B2(b[20]), .C1(n1), .C2(n1098), .A(n129), .ZN(
        n350) );
  INV_X2 U406 ( .A(n130), .ZN(\intadd_34/B[2] ) );
  INV_X2 U407 ( .A(\intadd_6/SUM[0] ), .ZN(\intadd_34/A[2] ) );
  NOR2_X1 U408 ( .A1(n654), .A2(n689), .ZN(n132) );
  AOI22_X1 U409 ( .A1(b[19]), .A2(n694), .B1(n693), .B2(n1106), .ZN(n131) );
  OAI221_X1 U410 ( .B1(b[18]), .B2(n690), .C1(n1114), .C2(n691), .A(n131), 
        .ZN(n838) );
  AOI21_X1 U411 ( .B1(n654), .B2(n689), .A(n1105), .ZN(n836) );
  OAI21_X1 U412 ( .B1(n132), .B2(n838), .A(n836), .ZN(n803) );
  AOI22_X1 U413 ( .A1(b[18]), .A2(n826), .B1(n825), .B2(n1114), .ZN(n133) );
  AOI221_X1 U414 ( .B1(n846), .B2(b[17]), .C1(n828), .C2(n824), .A(n133), .ZN(
        n802) );
  AOI22_X1 U415 ( .A1(b[15]), .A2(n884), .B1(n885), .B2(n687), .ZN(n134) );
  AOI221_X1 U416 ( .B1(n882), .B2(b[16]), .C1(n881), .C2(n575), .A(n134), .ZN(
        n801) );
  INV_X2 U417 ( .A(n135), .ZN(n152) );
  AOI22_X1 U418 ( .A1(b[20]), .A2(n813), .B1(n812), .B2(n1098), .ZN(n136) );
  AOI221_X1 U419 ( .B1(n816), .B2(b[19]), .C1(n815), .C2(n1106), .A(n136), 
        .ZN(n751) );
  AOI22_X1 U420 ( .A1(b[17]), .A2(n691), .B1(n690), .B2(n824), .ZN(n137) );
  AOI221_X1 U421 ( .B1(n694), .B2(b[18]), .C1(n693), .C2(n1114), .A(n137), 
        .ZN(n750) );
  NAND2_X1 U422 ( .A1(a[21]), .A2(a[22]), .ZN(n1164) );
  OAI21_X1 U423 ( .B1(a[21]), .B2(a[22]), .A(n1164), .ZN(n576) );
  NOR2_X1 U424 ( .A1(a[23]), .A2(n576), .ZN(n1139) );
  NOR2_X1 U425 ( .A1(n1105), .A2(n576), .ZN(n1147) );
  NAND2_X1 U426 ( .A1(n1162), .A2(n1105), .ZN(n1150) );
  NOR3_X1 U427 ( .A1(a[21]), .A2(a[22]), .A3(n1105), .ZN(n1141) );
  AOI22_X1 U428 ( .A1(b[9]), .A2(n1150), .B1(n1108), .B2(n689), .ZN(n138) );
  AOI221_X1 U429 ( .B1(n1139), .B2(b[10]), .C1(n1147), .C2(n649), .A(n138), 
        .ZN(n749) );
  NOR2_X1 U430 ( .A1(n1105), .A2(n654), .ZN(n747) );
  NOR2_X1 U431 ( .A1(a[8]), .A2(n767), .ZN(n139) );
  AOI221_X1 U432 ( .B1(n771), .B2(b[23]), .C1(n139), .C2(n1163), .A(n784), 
        .ZN(n748) );
  INV_X1 U433 ( .A(n748), .ZN(n143) );
  AOI22_X1 U434 ( .A1(b[22]), .A2(n791), .B1(n790), .B2(n1140), .ZN(n140) );
  AOI221_X1 U435 ( .B1(n819), .B2(b[21]), .C1(n793), .C2(n878), .A(n140), .ZN(
        n746) );
  OAI21_X1 U436 ( .B1(n748), .B2(n747), .A(n746), .ZN(n142) );
  AOI22_X1 U437 ( .A1(b[20]), .A2(n816), .B1(n815), .B2(n1098), .ZN(n141) );
  OAI221_X1 U438 ( .B1(b[21]), .B2(n812), .C1(n878), .C2(n813), .A(n141), .ZN(
        n145) );
  OAI211_X1 U439 ( .C1(n144), .C2(n143), .A(n142), .B(n145), .ZN(n796) );
  NAND2_X1 U440 ( .A1(n147), .A2(n146), .ZN(n795) );
  AOI21_X1 U441 ( .B1(n798), .B2(n796), .A(n148), .ZN(n151) );
  INV_X2 U442 ( .A(\intadd_14/SUM[0] ), .ZN(n150) );
  INV_X2 U443 ( .A(n149), .ZN(\intadd_1/B[4] ) );
  FA_X1 U444 ( .A(n152), .B(n151), .CI(n150), .CO(n153), .S(n149) );
  AOI22_X1 U445 ( .A1(b[20]), .A2(n884), .B1(n885), .B2(n1098), .ZN(n154) );
  AOI221_X1 U446 ( .B1(n882), .B2(b[21]), .C1(n881), .C2(n878), .A(n154), .ZN(
        n227) );
  NAND2_X1 U447 ( .A1(b[15]), .A2(b[14]), .ZN(n155) );
  OAI21_X1 U448 ( .B1(b[15]), .B2(b[14]), .A(a[23]), .ZN(n226) );
  AOI21_X1 U449 ( .B1(n227), .B2(n155), .A(n226), .ZN(n162) );
  OR3_X1 U450 ( .A1(a[19]), .A2(a[20]), .A3(n1095), .ZN(n623) );
  NOR2_X1 U451 ( .A1(n842), .A2(n156), .ZN(n289) );
  NAND2_X1 U452 ( .A1(n1095), .A2(n289), .ZN(n624) );
  OAI22_X1 U453 ( .A1(n842), .A2(n156), .B1(a[20]), .B2(a[19]), .ZN(n294) );
  NOR2_X1 U454 ( .A1(n294), .A2(a[21]), .ZN(n626) );
  NOR2_X1 U455 ( .A1(n294), .A2(n1095), .ZN(n1096) );
  AOI22_X1 U456 ( .A1(b[20]), .A2(n626), .B1(n1096), .B2(n1098), .ZN(n157) );
  OAI221_X1 U457 ( .B1(b[19]), .B2(n623), .C1(n1106), .C2(n624), .A(n157), 
        .ZN(n161) );
  AOI22_X1 U458 ( .A1(b[18]), .A2(n1139), .B1(n1147), .B2(n1114), .ZN(n158) );
  OAI221_X1 U459 ( .B1(b[17]), .B2(n1108), .C1(n824), .C2(n1150), .A(n158), 
        .ZN(n160) );
  INV_X1 U460 ( .A(n159), .ZN(\intadd_22/A[3] ) );
  FA_X1 U461 ( .A(n162), .B(n161), .CI(n160), .CO(n159), .S(n163) );
  INV_X1 U462 ( .A(n163), .ZN(\intadd_23/A[3] ) );
  FA_X1 U463 ( .A(n166), .B(n165), .CI(n164), .CO(n185), .S(n29) );
  NAND2_X1 U464 ( .A1(n784), .A2(n628), .ZN(n181) );
  AOI21_X1 U465 ( .B1(n769), .B2(n181), .A(b[0]), .ZN(n171) );
  XOR2_X1 U466 ( .A(n170), .B(n167), .Z(n174) );
  NAND2_X1 U467 ( .A1(n173), .A2(n168), .ZN(n169) );
  OAI211_X1 U468 ( .C1(n173), .C2(n170), .A(n171), .B(n169), .ZN(n184) );
  AOI21_X1 U469 ( .B1(n174), .B2(n173), .A(n171), .ZN(n172) );
  OAI21_X1 U470 ( .B1(n174), .B2(n173), .A(n172), .ZN(n182) );
  NAND2_X1 U471 ( .A1(n184), .A2(n182), .ZN(n175) );
  XNOR2_X1 U472 ( .A(n185), .B(n175), .ZN(n205) );
  AOI22_X1 U473 ( .A1(b[1]), .A2(n776), .B1(n725), .B2(n628), .ZN(n176) );
  OAI221_X1 U474 ( .B1(b[2]), .B2(n773), .C1(n606), .C2(n723), .A(n176), .ZN(
        n191) );
  NOR2_X1 U475 ( .A1(n1247), .A2(n768), .ZN(n190) );
  AOI22_X1 U476 ( .A1(b[3]), .A2(n729), .B1(n717), .B2(n555), .ZN(n177) );
  OAI221_X1 U477 ( .B1(b[4]), .B2(n714), .C1(n704), .C2(n715), .A(n177), .ZN(
        n189) );
  OAI221_X1 U478 ( .B1(a[1]), .B2(b[9]), .C1(n1239), .C2(n689), .A(a[0]), .ZN(
        n178) );
  OAI21_X1 U479 ( .B1(b[8]), .B2(n508), .A(n178), .ZN(n510) );
  NOR2_X1 U480 ( .A1(n771), .A2(n722), .ZN(n782) );
  OAI211_X1 U481 ( .C1(n1238), .C2(n767), .A(b[1]), .B(n179), .ZN(n180) );
  OAI221_X1 U482 ( .B1(n1238), .B2(n782), .C1(n1238), .C2(n181), .A(n180), 
        .ZN(n509) );
  AOI222_X1 U483 ( .A1(\intadd_0/SUM[0] ), .A2(n205), .B1(\intadd_0/SUM[0] ), 
        .B2(n204), .C1(n205), .C2(n204), .ZN(n216) );
  AOI21_X1 U484 ( .B1(n185), .B2(n184), .A(n183), .ZN(n543) );
  XOR2_X1 U485 ( .A(n216), .B(n218), .Z(n212) );
  INV_X2 U486 ( .A(\intadd_8/SUM[0] ), .ZN(n194) );
  FA_X1 U487 ( .A(n188), .B(n187), .CI(n186), .CO(n200), .S(n197) );
  FA_X1 U488 ( .A(n191), .B(n190), .CI(n189), .CO(n511), .S(n192) );
  NOR2_X1 U489 ( .A1(\intadd_8/SUM[1] ), .A2(n1053), .ZN(n1052) );
  FA_X1 U490 ( .A(n194), .B(n200), .CI(n201), .CO(n193), .S(n199) );
  FA_X1 U491 ( .A(n197), .B(n196), .CI(n195), .CO(n198), .S(n25) );
  NAND2_X1 U492 ( .A1(n199), .A2(n198), .ZN(n1051) );
  NAND2_X1 U493 ( .A1(\intadd_26/n1 ), .A2(n1051), .ZN(n1055) );
  NOR2_X1 U494 ( .A1(n199), .A2(n198), .ZN(n1050) );
  OAI21_X1 U495 ( .B1(n1050), .B2(n1053), .A(\intadd_8/SUM[1] ), .ZN(n203) );
  OR3_X1 U496 ( .A1(n1054), .A2(n201), .A3(n200), .ZN(n202) );
  OAI211_X1 U497 ( .C1(n1052), .C2(n1055), .A(n203), .B(n202), .ZN(n214) );
  AOI22_X1 U498 ( .A1(n207), .A2(n206), .B1(n205), .B2(n204), .ZN(n208) );
  XNOR2_X1 U499 ( .A(\intadd_0/SUM[0] ), .B(n208), .ZN(n213) );
  NAND2_X1 U500 ( .A1(n214), .A2(n213), .ZN(n211) );
  NAND2_X1 U501 ( .A1(n214), .A2(\intadd_8/n4 ), .ZN(n210) );
  NAND2_X1 U502 ( .A1(n213), .A2(\intadd_8/n4 ), .ZN(n209) );
  NAND3_X1 U503 ( .A1(n211), .A2(n210), .A3(n209), .ZN(n217) );
  XNOR2_X1 U504 ( .A(n212), .B(n217), .ZN(\d[11]_BAR ) );
  XOR2_X1 U505 ( .A(n214), .B(n213), .Z(n215) );
  XNOR2_X1 U506 ( .A(n215), .B(\intadd_8/n4 ), .ZN(\d[10]_BAR ) );
  NAND2_X1 U507 ( .A1(n216), .A2(n218), .ZN(n221) );
  NAND2_X1 U508 ( .A1(n216), .A2(n217), .ZN(n220) );
  NAND2_X1 U509 ( .A1(n218), .A2(n217), .ZN(n219) );
  NAND3_X1 U510 ( .A1(n221), .A2(n220), .A3(n219), .ZN(\intadd_8/n2 ) );
  AOI22_X1 U511 ( .A1(b[22]), .A2(n691), .B1(n690), .B2(n1140), .ZN(n222) );
  AOI221_X1 U512 ( .B1(n694), .B2(b[23]), .C1(n693), .C2(n1163), .A(n222), 
        .ZN(\intadd_23/B[0] ) );
  AOI22_X1 U513 ( .A1(b[18]), .A2(n884), .B1(n885), .B2(n1114), .ZN(n223) );
  AOI221_X1 U514 ( .B1(n882), .B2(b[19]), .C1(n881), .C2(n1106), .A(n223), 
        .ZN(\intadd_23/CI ) );
  NOR2_X1 U515 ( .A1(n637), .A2(n650), .ZN(n225) );
  AOI22_X1 U516 ( .A1(b[20]), .A2(n846), .B1(n828), .B2(n1098), .ZN(n224) );
  OAI221_X1 U517 ( .B1(b[21]), .B2(n825), .C1(n878), .C2(n826), .A(n224), .ZN(
        n244) );
  AOI21_X1 U518 ( .B1(n637), .B2(n650), .A(n1105), .ZN(n242) );
  OAI21_X1 U519 ( .B1(n225), .B2(n244), .A(n242), .ZN(\intadd_23/B[1] ) );
  AOI21_X1 U520 ( .B1(b[14]), .B2(b[15]), .A(n226), .ZN(n228) );
  XOR2_X1 U521 ( .A(n228), .B(n227), .Z(\intadd_23/B[2] ) );
  AOI22_X1 U522 ( .A1(b[15]), .A2(n1150), .B1(n1108), .B2(n687), .ZN(n229) );
  AOI221_X1 U523 ( .B1(n1139), .B2(b[16]), .C1(n1147), .C2(n575), .A(n229), 
        .ZN(\intadd_22/A[0] ) );
  AOI22_X1 U524 ( .A1(b[18]), .A2(n1103), .B1(n1104), .B2(n1114), .ZN(n230) );
  AOI221_X1 U525 ( .B1(n1101), .B2(b[17]), .C1(n1100), .C2(n824), .A(n230), 
        .ZN(\intadd_22/B[0] ) );
  AOI22_X1 U526 ( .A1(b[19]), .A2(n884), .B1(n885), .B2(n1106), .ZN(n231) );
  AOI221_X1 U527 ( .B1(n882), .B2(b[20]), .C1(n881), .C2(n1098), .A(n231), 
        .ZN(\intadd_22/CI ) );
  AOI22_X1 U528 ( .A1(b[23]), .A2(n826), .B1(n825), .B2(n1151), .ZN(n232) );
  AOI221_X1 U529 ( .B1(n846), .B2(b[22]), .C1(n828), .C2(n1140), .A(n232), 
        .ZN(\intadd_22/A[1] ) );
  NOR2_X1 U530 ( .A1(n1105), .A2(n554), .ZN(n238) );
  AOI22_X1 U531 ( .A1(b[22]), .A2(n826), .B1(n825), .B2(n1140), .ZN(n233) );
  AOI221_X1 U532 ( .B1(n846), .B2(b[21]), .C1(n828), .C2(n878), .A(n233), .ZN(
        n237) );
  AOI221_X1 U533 ( .B1(n235), .B2(b[23]), .C1(n234), .C2(n1163), .A(n693), 
        .ZN(n236) );
  FA_X1 U534 ( .A(n238), .B(n237), .CI(n236), .CO(\intadd_22/B[1] ), .S(
        \intadd_23/A[1] ) );
  AOI22_X1 U535 ( .A1(b[20]), .A2(n826), .B1(n825), .B2(n1098), .ZN(n239) );
  AOI221_X1 U536 ( .B1(n846), .B2(b[19]), .C1(n828), .C2(n1106), .A(n239), 
        .ZN(\intadd_35/A[0] ) );
  AOI22_X1 U537 ( .A1(b[17]), .A2(n884), .B1(n885), .B2(n824), .ZN(n240) );
  AOI221_X1 U538 ( .B1(n882), .B2(b[18]), .C1(n881), .C2(n1114), .A(n240), 
        .ZN(\intadd_35/B[0] ) );
  AOI22_X1 U539 ( .A1(b[13]), .A2(n1150), .B1(n1108), .B2(n637), .ZN(n241) );
  AOI221_X1 U540 ( .B1(n1147), .B2(n554), .C1(n1139), .C2(b[14]), .A(n241), 
        .ZN(\intadd_35/CI ) );
  OAI21_X1 U541 ( .B1(n637), .B2(n650), .A(n242), .ZN(n243) );
  XOR2_X1 U542 ( .A(n244), .B(n243), .Z(\intadd_35/B[1] ) );
  NOR2_X1 U543 ( .A1(a[12]), .A2(n245), .ZN(n247) );
  AOI221_X1 U544 ( .B1(n816), .B2(b[23]), .C1(n247), .C2(n1163), .A(n246), 
        .ZN(n256) );
  AOI22_X1 U545 ( .A1(b[21]), .A2(n691), .B1(n690), .B2(n878), .ZN(n248) );
  AOI221_X1 U546 ( .B1(n694), .B2(b[22]), .C1(n693), .C2(n1140), .A(n248), 
        .ZN(n255) );
  NOR2_X1 U547 ( .A1(n1105), .A2(n650), .ZN(n254) );
  AOI22_X1 U548 ( .A1(b[14]), .A2(n1150), .B1(n1108), .B2(n554), .ZN(n249) );
  AOI221_X1 U549 ( .B1(n1139), .B2(b[15]), .C1(n1147), .C2(n687), .A(n249), 
        .ZN(n264) );
  AOI22_X1 U550 ( .A1(b[17]), .A2(n1103), .B1(n1104), .B2(n824), .ZN(n250) );
  AOI221_X1 U551 ( .B1(n1101), .B2(b[16]), .C1(n1100), .C2(n575), .A(n250), 
        .ZN(n263) );
  AOI22_X1 U552 ( .A1(b[20]), .A2(n691), .B1(n690), .B2(n1098), .ZN(n251) );
  AOI221_X1 U553 ( .B1(n694), .B2(b[21]), .C1(n693), .C2(n878), .A(n251), .ZN(
        n806) );
  AOI22_X1 U554 ( .A1(b[15]), .A2(n1103), .B1(n1104), .B2(n687), .ZN(n252) );
  AOI221_X1 U555 ( .B1(n1101), .B2(b[14]), .C1(n1100), .C2(n554), .A(n252), 
        .ZN(n805) );
  AOI22_X1 U556 ( .A1(b[12]), .A2(n1150), .B1(n1108), .B2(n650), .ZN(n253) );
  AOI221_X1 U557 ( .B1(n1147), .B2(n637), .C1(n1139), .C2(b[13]), .A(n253), 
        .ZN(n804) );
  FA_X1 U558 ( .A(n256), .B(n255), .CI(n254), .CO(n265), .S(n799) );
  AOI22_X1 U559 ( .A1(b[19]), .A2(n826), .B1(n825), .B2(n1106), .ZN(n257) );
  AOI221_X1 U560 ( .B1(n846), .B2(b[18]), .C1(n828), .C2(n1114), .A(n257), 
        .ZN(n278) );
  NAND2_X1 U561 ( .A1(b[10]), .A2(b[11]), .ZN(n258) );
  OAI21_X1 U562 ( .B1(b[10]), .B2(b[11]), .A(a[23]), .ZN(n277) );
  AOI21_X1 U563 ( .B1(n278), .B2(n258), .A(n277), .ZN(n268) );
  AOI22_X1 U564 ( .A1(b[15]), .A2(n1101), .B1(n1100), .B2(n687), .ZN(n259) );
  OAI221_X1 U565 ( .B1(b[16]), .B2(n1104), .C1(n575), .C2(n1103), .A(n259), 
        .ZN(n267) );
  AOI22_X1 U566 ( .A1(b[23]), .A2(n813), .B1(n812), .B2(n1151), .ZN(n261) );
  AOI221_X1 U567 ( .B1(n816), .B2(b[22]), .C1(n815), .C2(n1140), .A(n261), 
        .ZN(n808) );
  AOI22_X1 U568 ( .A1(b[16]), .A2(n884), .B1(n885), .B2(n575), .ZN(n262) );
  AOI221_X1 U569 ( .B1(n882), .B2(b[17]), .C1(n881), .C2(n824), .A(n262), .ZN(
        n807) );
  INV_X1 U570 ( .A(n282), .ZN(n270) );
  FA_X1 U571 ( .A(n265), .B(n264), .CI(n263), .CO(\intadd_35/B[2] ), .S(n266)
         );
  INV_X1 U572 ( .A(n266), .ZN(n269) );
  NAND2_X1 U573 ( .A1(n268), .A2(n267), .ZN(n280) );
  INV_X1 U574 ( .A(n280), .ZN(n271) );
  AOI211_X1 U575 ( .C1(n281), .C2(n270), .A(n269), .B(n271), .ZN(n887) );
  INV_X1 U576 ( .A(n887), .ZN(n272) );
  OAI211_X1 U577 ( .C1(n271), .C2(n270), .A(n269), .B(n281), .ZN(n888) );
  NAND2_X1 U578 ( .A1(n272), .A2(n888), .ZN(n273) );
  XNOR2_X1 U579 ( .A(n889), .B(n273), .ZN(\intadd_14/A[3] ) );
  AOI22_X1 U580 ( .A1(b[14]), .A2(n1103), .B1(n1104), .B2(n554), .ZN(n274) );
  AOI221_X1 U581 ( .B1(n1101), .B2(b[13]), .C1(n1100), .C2(n637), .A(n274), 
        .ZN(\intadd_14/A[0] ) );
  AOI22_X1 U582 ( .A1(b[11]), .A2(n1150), .B1(n1108), .B2(n754), .ZN(n275) );
  AOI221_X1 U583 ( .B1(n1147), .B2(n650), .C1(n1139), .C2(b[12]), .A(n275), 
        .ZN(\intadd_14/B[0] ) );
  AOI22_X1 U584 ( .A1(b[19]), .A2(n691), .B1(n690), .B2(n1106), .ZN(n276) );
  AOI221_X1 U585 ( .B1(n694), .B2(b[20]), .C1(n693), .C2(n1098), .A(n276), 
        .ZN(\intadd_14/CI ) );
  AOI21_X1 U586 ( .B1(b[11]), .B2(b[10]), .A(n277), .ZN(n279) );
  XOR2_X1 U587 ( .A(n279), .B(n278), .Z(\intadd_14/B[1] ) );
  NAND2_X1 U588 ( .A1(n281), .A2(n280), .ZN(n283) );
  XNOR2_X1 U589 ( .A(n283), .B(n282), .ZN(\intadd_14/B[2] ) );
  AOI22_X1 U590 ( .A1(b[19]), .A2(n1103), .B1(n1104), .B2(n1106), .ZN(n284) );
  AOI221_X1 U591 ( .B1(n1101), .B2(b[18]), .C1(n1100), .C2(n1114), .A(n284), 
        .ZN(n287) );
  AOI22_X1 U592 ( .A1(b[16]), .A2(n1150), .B1(n1108), .B2(n575), .ZN(n285) );
  AOI221_X1 U593 ( .B1(n1147), .B2(n824), .C1(n1139), .C2(b[17]), .A(n285), 
        .ZN(n286) );
  FA_X1 U594 ( .A(n288), .B(n287), .CI(n286), .CO(\intadd_22/B[2] ), .S(
        \intadd_23/A[2] ) );
  NOR2_X1 U595 ( .A1(n289), .A2(n1095), .ZN(n1161) );
  NAND2_X1 U596 ( .A1(n1161), .A2(n1238), .ZN(n290) );
  AOI21_X1 U597 ( .B1(b[1]), .B2(n623), .A(n290), .ZN(n337) );
  OAI211_X1 U598 ( .C1(n624), .C2(n1238), .A(n623), .B(n290), .ZN(n291) );
  AOI221_X1 U599 ( .B1(n626), .B2(b[1]), .C1(n1096), .C2(n628), .A(n291), .ZN(
        n292) );
  NOR2_X1 U600 ( .A1(n337), .A2(n292), .ZN(\intadd_34/A[1] ) );
  AOI22_X1 U601 ( .A1(b[2]), .A2(n882), .B1(n881), .B2(n606), .ZN(n293) );
  OAI221_X1 U602 ( .B1(b[1]), .B2(n885), .C1(n628), .C2(n884), .A(n293), .ZN(
        \intadd_34/A[0] ) );
  NOR2_X1 U603 ( .A1(n294), .A2(n1247), .ZN(\intadd_34/B[0] ) );
  AOI22_X1 U604 ( .A1(b[3]), .A2(n846), .B1(n828), .B2(n555), .ZN(n295) );
  OAI221_X1 U605 ( .B1(b[4]), .B2(n825), .C1(n704), .C2(n826), .A(n295), .ZN(
        \intadd_34/CI ) );
  AOI22_X1 U606 ( .A1(b[8]), .A2(n816), .B1(n815), .B2(n654), .ZN(n296) );
  OAI221_X1 U607 ( .B1(b[9]), .B2(n812), .C1(n689), .C2(n813), .A(n296), .ZN(
        \intadd_34/B[1] ) );
  AOI22_X1 U608 ( .A1(b[22]), .A2(n528), .B1(n527), .B2(n1140), .ZN(n297) );
  AOI21_X1 U609 ( .B1(n530), .B2(n878), .A(n297), .ZN(\intadd_6/A[0] ) );
  AOI22_X1 U610 ( .A1(b[6]), .A2(n826), .B1(n825), .B2(n764), .ZN(n298) );
  AOI221_X1 U611 ( .B1(n846), .B2(b[5]), .C1(n828), .C2(n741), .A(n298), .ZN(
        \intadd_6/B[0] ) );
  AOI22_X1 U612 ( .A1(b[7]), .A2(n691), .B1(n690), .B2(n712), .ZN(n299) );
  AOI221_X1 U613 ( .B1(n694), .B2(b[8]), .C1(n693), .C2(n654), .A(n299), .ZN(
        \intadd_6/CI ) );
  AOI22_X1 U614 ( .A1(b[3]), .A2(n826), .B1(n825), .B2(n555), .ZN(n300) );
  AOI221_X1 U615 ( .B1(n846), .B2(b[2]), .C1(n828), .C2(n606), .A(n300), .ZN(
        n405) );
  AOI22_X1 U616 ( .A1(b[11]), .A2(n780), .B1(n720), .B2(n754), .ZN(n301) );
  AOI221_X1 U617 ( .B1(n771), .B2(b[10]), .C1(n722), .C2(n649), .A(n301), .ZN(
        n404) );
  AOI22_X1 U618 ( .A1(b[4]), .A2(n691), .B1(n690), .B2(n704), .ZN(n302) );
  AOI221_X1 U619 ( .B1(n694), .B2(b[5]), .C1(n693), .C2(n741), .A(n302), .ZN(
        n403) );
  AOI22_X1 U620 ( .A1(b[7]), .A2(n813), .B1(n812), .B2(n712), .ZN(n303) );
  AOI221_X1 U621 ( .B1(n816), .B2(b[6]), .C1(n815), .C2(n764), .A(n303), .ZN(
        n311) );
  AOI22_X1 U622 ( .A1(b[19]), .A2(n528), .B1(n527), .B2(n1106), .ZN(n304) );
  AOI21_X1 U623 ( .B1(n530), .B2(n1114), .A(n304), .ZN(n310) );
  NOR2_X1 U624 ( .A1(n311), .A2(n310), .ZN(n409) );
  OAI21_X1 U625 ( .B1(n776), .B2(n725), .A(n305), .ZN(n306) );
  OAI221_X1 U626 ( .B1(b[13]), .B2(n773), .C1(n637), .C2(n723), .A(n306), .ZN(
        n411) );
  AOI22_X1 U627 ( .A1(b[15]), .A2(n715), .B1(n714), .B2(n687), .ZN(n307) );
  AOI221_X1 U628 ( .B1(n729), .B2(b[14]), .C1(n717), .C2(n554), .A(n307), .ZN(
        n418) );
  AOI22_X1 U629 ( .A1(b[17]), .A2(n633), .B1(n1), .B2(n824), .ZN(n308) );
  OAI221_X1 U630 ( .B1(b[16]), .B2(n631), .C1(n575), .C2(n643), .A(n308), .ZN(
        n313) );
  AOI22_X1 U631 ( .A1(b[8]), .A2(n819), .B1(n793), .B2(n654), .ZN(n309) );
  OAI221_X1 U632 ( .B1(b[9]), .B2(n790), .C1(n689), .C2(n791), .A(n309), .ZN(
        n312) );
  NAND2_X1 U633 ( .A1(n313), .A2(n312), .ZN(n416) );
  NAND2_X1 U634 ( .A1(n311), .A2(n310), .ZN(n317) );
  NOR2_X1 U635 ( .A1(n313), .A2(n312), .ZN(n315) );
  AOI211_X1 U636 ( .C1(n418), .C2(n416), .A(n410), .B(n315), .ZN(n314) );
  OAI21_X1 U637 ( .B1(n409), .B2(n411), .A(n314), .ZN(n399) );
  INV_X1 U638 ( .A(n418), .ZN(n316) );
  AOI22_X1 U639 ( .A1(n411), .A2(n317), .B1(n316), .B2(n417), .ZN(n319) );
  NAND3_X1 U640 ( .A1(n319), .A2(n318), .A3(n416), .ZN(n400) );
  AOI21_X1 U641 ( .B1(n401), .B2(n399), .A(n320), .ZN(\intadd_32/A[1] ) );
  AOI22_X1 U642 ( .A1(b[12]), .A2(n780), .B1(n720), .B2(n650), .ZN(n321) );
  AOI221_X1 U643 ( .B1(n771), .B2(b[11]), .C1(n722), .C2(n754), .A(n321), .ZN(
        \intadd_33/A[0] ) );
  AOI22_X1 U644 ( .A1(b[10]), .A2(n791), .B1(n790), .B2(n649), .ZN(n322) );
  AOI221_X1 U645 ( .B1(n819), .B2(b[9]), .C1(n793), .C2(n689), .A(n322), .ZN(
        \intadd_33/B[0] ) );
  AOI22_X1 U646 ( .A1(b[17]), .A2(n643), .B1(n631), .B2(n824), .ZN(n323) );
  AOI221_X1 U647 ( .B1(n633), .B2(b[18]), .C1(n1), .C2(n1114), .A(n323), .ZN(
        \intadd_33/CI ) );
  AOI22_X1 U648 ( .A1(b[13]), .A2(n780), .B1(n720), .B2(n637), .ZN(n324) );
  AOI221_X1 U649 ( .B1(n771), .B2(b[12]), .C1(n722), .C2(n650), .A(n324), .ZN(
        \intadd_7/A[0] ) );
  AOI22_X1 U650 ( .A1(b[5]), .A2(n826), .B1(n825), .B2(n741), .ZN(n325) );
  AOI221_X1 U651 ( .B1(n846), .B2(b[4]), .C1(n828), .C2(n704), .A(n325), .ZN(
        \intadd_7/B[0] ) );
  AOI22_X1 U652 ( .A1(b[2]), .A2(n884), .B1(n885), .B2(n606), .ZN(n326) );
  AOI221_X1 U653 ( .B1(n882), .B2(b[3]), .C1(n881), .C2(n555), .A(n326), .ZN(
        \intadd_7/CI ) );
  NAND2_X1 U654 ( .A1(b[0]), .A2(n701), .ZN(\intadd_24/A[0] ) );
  AOI22_X1 U655 ( .A1(b[1]), .A2(n624), .B1(n623), .B2(n628), .ZN(n327) );
  AOI221_X1 U656 ( .B1(n626), .B2(b[2]), .C1(n1096), .C2(n606), .A(n327), .ZN(
        \intadd_24/B[0] ) );
  AOI22_X1 U657 ( .A1(b[3]), .A2(n884), .B1(n885), .B2(n555), .ZN(n328) );
  AOI221_X1 U658 ( .B1(n882), .B2(b[4]), .C1(n881), .C2(n704), .A(n328), .ZN(
        \intadd_24/CI ) );
  XNOR2_X1 U659 ( .A(n330), .B(n329), .ZN(\intadd_10/B[1] ) );
  AOI22_X1 U660 ( .A1(b[3]), .A2(n691), .B1(n690), .B2(n555), .ZN(n332) );
  AOI221_X1 U661 ( .B1(n694), .B2(b[4]), .C1(n693), .C2(n704), .A(n332), .ZN(
        \intadd_10/B[0] ) );
  AOI22_X1 U662 ( .A1(b[2]), .A2(n826), .B1(n825), .B2(n606), .ZN(n333) );
  AOI221_X1 U663 ( .B1(n846), .B2(b[1]), .C1(n828), .C2(n628), .A(n333), .ZN(
        \intadd_10/CI ) );
  FA_X1 U664 ( .A(n336), .B(n335), .CI(n334), .CO(\intadd_33/B[1] ), .S(n126)
         );
  AOI21_X1 U665 ( .B1(n342), .B2(n341), .A(n340), .ZN(n338) );
  OAI211_X1 U666 ( .C1(n342), .C2(n341), .A(n343), .B(n339), .ZN(n385) );
  FA_X1 U667 ( .A(n342), .B(n341), .CI(n340), .CO(n344), .S(n110) );
  NOR2_X1 U668 ( .A1(n344), .A2(n343), .ZN(n387) );
  NOR2_X1 U669 ( .A1(n345), .A2(n387), .ZN(n349) );
  FA_X1 U670 ( .A(n348), .B(n347), .CI(n346), .CO(n384), .S(n117) );
  XOR2_X1 U671 ( .A(n349), .B(n384), .Z(\intadd_33/B[2] ) );
  FA_X1 U672 ( .A(n352), .B(n351), .CI(n350), .CO(\intadd_24/A[1] ), .S(n130)
         );
  AOI22_X1 U673 ( .A1(b[16]), .A2(n723), .B1(n773), .B2(n575), .ZN(n353) );
  AOI221_X1 U674 ( .B1(n776), .B2(b[15]), .C1(n725), .C2(n687), .A(n353), .ZN(
        n361) );
  NAND2_X1 U675 ( .A1(n829), .A2(n554), .ZN(n355) );
  OAI22_X1 U676 ( .A1(n829), .A2(b[13]), .B1(n355), .B2(a[9]), .ZN(n354) );
  AOI21_X1 U677 ( .B1(n355), .B2(a[9]), .A(n354), .ZN(n357) );
  AOI22_X1 U678 ( .A1(n722), .A2(n637), .B1(n357), .B2(n356), .ZN(n360) );
  AOI22_X1 U679 ( .A1(b[18]), .A2(n715), .B1(n714), .B2(n1114), .ZN(n358) );
  AOI221_X1 U680 ( .B1(n729), .B2(b[17]), .C1(n717), .C2(n824), .A(n358), .ZN(
        n359) );
  FA_X1 U681 ( .A(n361), .B(n360), .CI(n359), .CO(\intadd_24/B[1] ), .S(
        \intadd_7/A[1] ) );
  AOI22_X1 U682 ( .A1(b[19]), .A2(n715), .B1(n714), .B2(n1106), .ZN(n362) );
  AOI221_X1 U683 ( .B1(n729), .B2(b[18]), .C1(n717), .C2(n1114), .A(n362), 
        .ZN(\intadd_16/A[0] ) );
  AOI22_X1 U684 ( .A1(b[7]), .A2(n826), .B1(n825), .B2(n712), .ZN(n363) );
  AOI221_X1 U685 ( .B1(n846), .B2(b[6]), .C1(n828), .C2(n764), .A(n363), .ZN(
        \intadd_16/B[0] ) );
  AOI22_X1 U686 ( .A1(b[8]), .A2(n691), .B1(n690), .B2(n654), .ZN(n364) );
  AOI221_X1 U687 ( .B1(n694), .B2(b[9]), .C1(n693), .C2(n689), .A(n364), .ZN(
        \intadd_16/CI ) );
  AOI22_X1 U688 ( .A1(b[15]), .A2(n780), .B1(n720), .B2(n687), .ZN(n365) );
  AOI221_X1 U689 ( .B1(n771), .B2(b[14]), .C1(n722), .C2(n554), .A(n365), .ZN(
        n390) );
  AOI22_X1 U690 ( .A1(b[17]), .A2(n723), .B1(n773), .B2(n824), .ZN(n366) );
  AOI221_X1 U691 ( .B1(n776), .B2(b[16]), .C1(n725), .C2(n575), .A(n366), .ZN(
        n389) );
  NOR2_X1 U692 ( .A1(n1141), .A2(n1138), .ZN(n605) );
  NAND2_X1 U693 ( .A1(a[23]), .A2(b[0]), .ZN(n636) );
  AOI221_X1 U694 ( .B1(b[1]), .B2(n367), .C1(n628), .C2(n636), .A(n576), .ZN(
        n368) );
  AOI21_X1 U695 ( .B1(b[0]), .B2(n369), .A(n368), .ZN(n388) );
  AOI22_X1 U696 ( .A1(b[8]), .A2(n826), .B1(n825), .B2(n654), .ZN(n370) );
  AOI221_X1 U697 ( .B1(n846), .B2(b[7]), .C1(n828), .C2(n712), .A(n370), .ZN(
        \intadd_27/A[0] ) );
  AOI22_X1 U698 ( .A1(b[20]), .A2(n715), .B1(n714), .B2(n1098), .ZN(n371) );
  AOI221_X1 U699 ( .B1(n729), .B2(b[19]), .C1(n717), .C2(n1106), .A(n371), 
        .ZN(\intadd_27/B[0] ) );
  AOI22_X1 U700 ( .A1(b[18]), .A2(n723), .B1(n773), .B2(n1114), .ZN(n372) );
  AOI221_X1 U701 ( .B1(n776), .B2(b[17]), .C1(n725), .C2(n824), .A(n372), .ZN(
        \intadd_27/CI ) );
  NOR2_X1 U702 ( .A1(n373), .A2(n878), .ZN(n375) );
  OAI22_X1 U703 ( .A1(n1098), .A2(n661), .B1(n375), .B2(a[3]), .ZN(n374) );
  AOI21_X1 U704 ( .B1(n375), .B2(a[3]), .A(n374), .ZN(n377) );
  AOI22_X1 U705 ( .A1(b[20]), .A2(n378), .B1(n377), .B2(n376), .ZN(n383) );
  AOI22_X1 U706 ( .A1(b[11]), .A2(n813), .B1(n812), .B2(n754), .ZN(n379) );
  AOI221_X1 U707 ( .B1(n816), .B2(b[10]), .C1(n815), .C2(n649), .A(n379), .ZN(
        n382) );
  AOI221_X1 U708 ( .B1(b[23]), .B2(a[1]), .C1(n1163), .C2(n1239), .A(n1246), 
        .ZN(n380) );
  AOI21_X1 U709 ( .B1(n530), .B2(n1140), .A(n380), .ZN(n381) );
  FA_X1 U710 ( .A(n383), .B(n382), .CI(n381), .CO(\intadd_16/A[1] ), .S(
        \intadd_6/B[1] ) );
  OAI21_X1 U711 ( .B1(n387), .B2(n386), .A(n385), .ZN(n396) );
  FA_X1 U712 ( .A(n390), .B(n389), .CI(n388), .CO(\intadd_24/A[2] ), .S(n395)
         );
  AOI22_X1 U713 ( .A1(b[4]), .A2(n884), .B1(n885), .B2(n704), .ZN(n391) );
  AOI221_X1 U714 ( .B1(n882), .B2(b[5]), .C1(n881), .C2(n741), .A(n391), .ZN(
        n612) );
  AOI22_X1 U715 ( .A1(b[3]), .A2(n1103), .B1(n1104), .B2(n555), .ZN(n392) );
  AOI221_X1 U716 ( .B1(n1101), .B2(b[2]), .C1(n1100), .C2(n606), .A(n392), 
        .ZN(n611) );
  AOI22_X1 U717 ( .A1(b[13]), .A2(n791), .B1(n790), .B2(n637), .ZN(n393) );
  AOI221_X1 U718 ( .B1(n819), .B2(b[12]), .C1(n793), .C2(n650), .A(n393), .ZN(
        n610) );
  FA_X1 U719 ( .A(n396), .B(n395), .CI(n394), .CO(\intadd_7/A[3] ), .S(n1001)
         );
  INV_X2 U720 ( .A(\intadd_32/n1 ), .ZN(n1000) );
  NAND2_X1 U721 ( .A1(n397), .A2(n1000), .ZN(n902) );
  NAND2_X1 U722 ( .A1(n902), .A2(n925), .ZN(n398) );
  XNOR2_X1 U723 ( .A(n398), .B(\intadd_7/SUM[2] ), .ZN(\intadd_11/B[3] ) );
  NAND2_X1 U724 ( .A1(n400), .A2(n399), .ZN(n402) );
  XNOR2_X1 U725 ( .A(n402), .B(n401), .ZN(\intadd_9/A[3] ) );
  FA_X1 U726 ( .A(n405), .B(n404), .CI(n403), .CO(n401), .S(\intadd_9/A[2] )
         );
  AOI22_X1 U727 ( .A1(b[2]), .A2(n691), .B1(n690), .B2(n606), .ZN(n406) );
  AOI221_X1 U728 ( .B1(n694), .B2(b[3]), .C1(n693), .C2(n555), .A(n406), .ZN(
        \intadd_9/A[0] ) );
  AOI22_X1 U729 ( .A1(b[7]), .A2(n791), .B1(n790), .B2(n712), .ZN(n407) );
  AOI221_X1 U730 ( .B1(n819), .B2(b[6]), .C1(n793), .C2(n764), .A(n407), .ZN(
        \intadd_9/B[0] ) );
  AOI22_X1 U731 ( .A1(b[5]), .A2(n813), .B1(n812), .B2(n741), .ZN(n408) );
  AOI221_X1 U732 ( .B1(n816), .B2(b[4]), .C1(n815), .C2(n704), .A(n408), .ZN(
        \intadd_9/CI ) );
  NOR2_X1 U733 ( .A1(n410), .A2(n409), .ZN(n412) );
  XNOR2_X1 U734 ( .A(n412), .B(n411), .ZN(n422) );
  AOI22_X1 U735 ( .A1(b[18]), .A2(n528), .B1(n527), .B2(n1114), .ZN(n413) );
  AOI21_X1 U736 ( .B1(n530), .B2(n824), .A(n413), .ZN(n428) );
  AOI22_X1 U737 ( .A1(b[8]), .A2(n791), .B1(n790), .B2(n654), .ZN(n414) );
  AOI221_X1 U738 ( .B1(n819), .B2(b[7]), .C1(n793), .C2(n712), .A(n414), .ZN(
        n427) );
  AOI22_X1 U739 ( .A1(b[6]), .A2(n813), .B1(n812), .B2(n764), .ZN(n415) );
  AOI221_X1 U740 ( .B1(n816), .B2(b[5]), .C1(n815), .C2(n741), .A(n415), .ZN(
        n426) );
  NAND2_X1 U741 ( .A1(n417), .A2(n416), .ZN(n419) );
  XNOR2_X1 U742 ( .A(n419), .B(n418), .ZN(n420) );
  FA_X1 U743 ( .A(n422), .B(n421), .CI(n420), .CO(\intadd_10/B[2] ), .S(
        \intadd_21/A[3] ) );
  AOI22_X1 U744 ( .A1(b[13]), .A2(n643), .B1(n631), .B2(n637), .ZN(n423) );
  AOI221_X1 U745 ( .B1(n633), .B2(b[14]), .C1(n1), .C2(n554), .A(n423), .ZN(
        \intadd_21/A[0] ) );
  AOI22_X1 U746 ( .A1(b[12]), .A2(n715), .B1(n714), .B2(n650), .ZN(n424) );
  AOI221_X1 U747 ( .B1(n729), .B2(b[11]), .C1(n717), .C2(n754), .A(n424), .ZN(
        \intadd_21/B[0] ) );
  AOI22_X1 U748 ( .A1(b[10]), .A2(n723), .B1(n773), .B2(n649), .ZN(n425) );
  AOI221_X1 U749 ( .B1(n776), .B2(b[9]), .C1(n725), .C2(n689), .A(n425), .ZN(
        \intadd_21/CI ) );
  FA_X1 U750 ( .A(n428), .B(n427), .CI(n426), .CO(n421), .S(\intadd_21/B[2] )
         );
  OAI22_X1 U751 ( .A1(b[8]), .A2(n769), .B1(n768), .B2(n429), .ZN(n430) );
  AOI21_X1 U752 ( .B1(n771), .B2(b[8]), .A(n430), .ZN(n439) );
  AOI221_X1 U753 ( .B1(a[1]), .B2(b[17]), .C1(n1239), .C2(n824), .A(n1246), 
        .ZN(n431) );
  AOI21_X1 U754 ( .B1(n530), .B2(n575), .A(n431), .ZN(n438) );
  AOI22_X1 U755 ( .A1(b[14]), .A2(n643), .B1(n631), .B2(n554), .ZN(n432) );
  AOI221_X1 U756 ( .B1(n633), .B2(b[15]), .C1(n1), .C2(n687), .A(n432), .ZN(
        n437) );
  AOI22_X1 U757 ( .A1(b[14]), .A2(n715), .B1(n714), .B2(n554), .ZN(n433) );
  AOI221_X1 U758 ( .B1(n729), .B2(b[13]), .C1(n717), .C2(n637), .A(n433), .ZN(
        n434) );
  FA_X1 U759 ( .A(n436), .B(n435), .CI(n434), .CO(\intadd_9/B[2] ), .S(
        \intadd_31/A[1] ) );
  FA_X1 U760 ( .A(n439), .B(n438), .CI(n437), .CO(n435), .S(\intadd_31/A[0] )
         );
  AOI22_X1 U761 ( .A1(b[3]), .A2(n813), .B1(n812), .B2(n555), .ZN(n440) );
  AOI221_X1 U762 ( .B1(n816), .B2(b[2]), .C1(n815), .C2(n606), .A(n440), .ZN(
        n465) );
  AOI22_X1 U763 ( .A1(b[5]), .A2(n791), .B1(n790), .B2(n741), .ZN(n441) );
  AOI221_X1 U764 ( .B1(n819), .B2(b[4]), .C1(n793), .C2(n704), .A(n441), .ZN(
        n464) );
  AOI22_X1 U765 ( .A1(b[9]), .A2(n723), .B1(n773), .B2(n689), .ZN(n442) );
  AOI221_X1 U766 ( .B1(n776), .B2(b[8]), .C1(n725), .C2(n654), .A(n442), .ZN(
        n463) );
  NOR2_X1 U767 ( .A1(n443), .A2(n449), .ZN(n470) );
  AOI22_X1 U768 ( .A1(b[11]), .A2(n715), .B1(n714), .B2(n754), .ZN(n444) );
  AOI221_X1 U769 ( .B1(n729), .B2(b[10]), .C1(n717), .C2(n649), .A(n444), .ZN(
        n468) );
  AOI22_X1 U770 ( .A1(b[15]), .A2(n528), .B1(n527), .B2(n687), .ZN(n445) );
  AOI21_X1 U771 ( .B1(n530), .B2(n554), .A(n445), .ZN(n467) );
  AOI22_X1 U772 ( .A1(b[7]), .A2(n780), .B1(n720), .B2(n712), .ZN(n446) );
  AOI221_X1 U773 ( .B1(n771), .B2(b[6]), .C1(n722), .C2(n764), .A(n446), .ZN(
        n466) );
  AOI21_X1 U774 ( .B1(n464), .B2(n463), .A(n465), .ZN(n447) );
  OAI211_X1 U775 ( .C1(n464), .C2(n463), .A(n449), .B(n448), .ZN(n469) );
  OAI21_X1 U776 ( .B1(n470), .B2(n450), .A(n469), .ZN(\intadd_31/B[0] ) );
  FA_X1 U777 ( .A(n453), .B(n452), .CI(n451), .CO(\intadd_21/B[1] ), .S(n70)
         );
  FA_X1 U778 ( .A(n456), .B(n455), .CI(n454), .CO(n88), .S(\intadd_30/B[0] )
         );
  FA_X1 U779 ( .A(n459), .B(n458), .CI(n457), .CO(\intadd_21/A[2] ), .S(n81)
         );
  AOI22_X1 U780 ( .A1(b[8]), .A2(n723), .B1(n773), .B2(n654), .ZN(n460) );
  AOI221_X1 U781 ( .B1(n776), .B2(b[7]), .C1(n725), .C2(n712), .A(n460), .ZN(
        \intadd_19/A[0] ) );
  AOI22_X1 U782 ( .A1(b[6]), .A2(n780), .B1(n720), .B2(n764), .ZN(n461) );
  AOI221_X1 U783 ( .B1(n771), .B2(b[5]), .C1(n722), .C2(n741), .A(n461), .ZN(
        \intadd_19/B[0] ) );
  AOI22_X1 U784 ( .A1(b[14]), .A2(n528), .B1(n527), .B2(n554), .ZN(n462) );
  AOI21_X1 U785 ( .B1(n530), .B2(n637), .A(n462), .ZN(\intadd_19/CI ) );
  FA_X1 U786 ( .A(n465), .B(n464), .CI(n463), .CO(n443), .S(\intadd_19/A[1] )
         );
  FA_X1 U787 ( .A(n468), .B(n467), .CI(n466), .CO(n472), .S(\intadd_19/B[1] )
         );
  NOR2_X1 U788 ( .A1(n471), .A2(n470), .ZN(n473) );
  XOR2_X1 U789 ( .A(n473), .B(n472), .Z(\intadd_19/B[2] ) );
  AOI22_X1 U790 ( .A1(b[5]), .A2(n780), .B1(n720), .B2(n741), .ZN(n474) );
  AOI221_X1 U791 ( .B1(n771), .B2(b[4]), .C1(n722), .C2(n704), .A(n474), .ZN(
        \intadd_20/A[0] ) );
  AOI22_X1 U792 ( .A1(b[9]), .A2(n715), .B1(n714), .B2(n689), .ZN(n475) );
  AOI221_X1 U793 ( .B1(n729), .B2(b[8]), .C1(n717), .C2(n654), .A(n475), .ZN(
        \intadd_20/B[0] ) );
  AOI22_X1 U794 ( .A1(b[3]), .A2(n791), .B1(n790), .B2(n555), .ZN(n476) );
  AOI221_X1 U795 ( .B1(n819), .B2(b[2]), .C1(n793), .C2(n606), .A(n476), .ZN(
        \intadd_20/CI ) );
  AOI22_X1 U796 ( .A1(b[11]), .A2(n528), .B1(n527), .B2(n754), .ZN(n477) );
  AOI21_X1 U797 ( .B1(n530), .B2(n649), .A(n477), .ZN(\intadd_18/A[0] ) );
  AOI22_X1 U798 ( .A1(b[7]), .A2(n715), .B1(n714), .B2(n712), .ZN(n478) );
  AOI221_X1 U799 ( .B1(n729), .B2(b[6]), .C1(n717), .C2(n764), .A(n478), .ZN(
        \intadd_18/B[0] ) );
  AOI22_X1 U800 ( .A1(b[3]), .A2(n780), .B1(n720), .B2(n555), .ZN(n479) );
  AOI221_X1 U801 ( .B1(n771), .B2(b[2]), .C1(n722), .C2(n606), .A(n479), .ZN(
        \intadd_18/CI ) );
  OAI222_X1 U802 ( .A1(b[0]), .A2(a[11]), .B1(n1238), .B2(n480), .C1(n819), 
        .C2(n793), .ZN(n481) );
  OAI221_X1 U803 ( .B1(b[1]), .B2(n790), .C1(n628), .C2(n791), .A(n481), .ZN(
        n499) );
  NAND3_X1 U804 ( .A1(n1238), .A2(n499), .A3(n818), .ZN(\intadd_18/A[1] ) );
  AOI22_X1 U805 ( .A1(b[9]), .A2(n643), .B1(n631), .B2(n689), .ZN(n482) );
  AOI221_X1 U806 ( .B1(n633), .B2(b[10]), .C1(n1), .C2(n649), .A(n482), .ZN(
        \intadd_18/B[1] ) );
  AOI22_X1 U807 ( .A1(b[10]), .A2(n643), .B1(n631), .B2(n649), .ZN(n483) );
  AOI221_X1 U808 ( .B1(n633), .B2(b[11]), .C1(n1), .C2(n754), .A(n483), .ZN(
        n488) );
  AOI22_X1 U809 ( .A1(b[7]), .A2(n723), .B1(n773), .B2(n712), .ZN(n484) );
  AOI221_X1 U810 ( .B1(n776), .B2(b[6]), .C1(n725), .C2(n764), .A(n484), .ZN(
        n487) );
  AOI221_X1 U811 ( .B1(a[1]), .B2(b[13]), .C1(n1239), .C2(n637), .A(n1246), 
        .ZN(n485) );
  AOI21_X1 U812 ( .B1(n530), .B2(n650), .A(n485), .ZN(n486) );
  FA_X1 U813 ( .A(n488), .B(n487), .CI(n486), .CO(\intadd_20/B[1] ), .S(
        \intadd_18/A[2] ) );
  XNOR2_X1 U814 ( .A(n490), .B(n489), .ZN(\intadd_29/A[1] ) );
  AOI22_X1 U815 ( .A1(b[8]), .A2(n715), .B1(n714), .B2(n654), .ZN(n491) );
  AOI221_X1 U816 ( .B1(n729), .B2(b[7]), .C1(n717), .C2(n712), .A(n491), .ZN(
        \intadd_29/A[0] ) );
  AOI22_X1 U817 ( .A1(b[6]), .A2(n723), .B1(n773), .B2(n764), .ZN(n492) );
  AOI221_X1 U818 ( .B1(n776), .B2(b[5]), .C1(n725), .C2(n741), .A(n492), .ZN(
        \intadd_29/B[0] ) );
  AOI221_X1 U819 ( .B1(a[1]), .B2(b[12]), .C1(n1239), .C2(n650), .A(n1246), 
        .ZN(n493) );
  AOI21_X1 U820 ( .B1(n530), .B2(n754), .A(n493), .ZN(\intadd_29/CI ) );
  FA_X1 U821 ( .A(n496), .B(n495), .CI(n494), .CO(n54), .S(\intadd_28/A[1] )
         );
  OAI21_X1 U822 ( .B1(n497), .B2(n1247), .A(n818), .ZN(n498) );
  XNOR2_X1 U823 ( .A(n499), .B(n498), .ZN(\intadd_28/A[0] ) );
  AOI22_X1 U824 ( .A1(b[4]), .A2(n776), .B1(n725), .B2(n704), .ZN(n500) );
  OAI221_X1 U825 ( .B1(b[5]), .B2(n773), .C1(n741), .C2(n723), .A(n500), .ZN(
        \intadd_28/B[0] ) );
  AOI22_X1 U826 ( .A1(b[9]), .A2(n633), .B1(n1), .B2(n689), .ZN(n501) );
  OAI221_X1 U827 ( .B1(b[8]), .B2(n631), .C1(n654), .C2(n643), .A(n501), .ZN(
        \intadd_28/CI ) );
  AOI22_X1 U828 ( .A1(b[7]), .A2(n643), .B1(n631), .B2(n712), .ZN(n502) );
  AOI221_X1 U829 ( .B1(n633), .B2(b[8]), .C1(n1), .C2(n654), .A(n502), .ZN(
        \intadd_0/A[0] ) );
  AOI22_X1 U830 ( .A1(b[6]), .A2(n715), .B1(n714), .B2(n764), .ZN(n503) );
  AOI221_X1 U831 ( .B1(n729), .B2(b[5]), .C1(n717), .C2(n741), .A(n503), .ZN(
        \intadd_0/B[0] ) );
  AOI22_X1 U832 ( .A1(b[10]), .A2(n528), .B1(n527), .B2(n649), .ZN(n504) );
  AOI21_X1 U833 ( .B1(n530), .B2(n689), .A(n504), .ZN(\intadd_0/CI ) );
  NOR2_X1 U834 ( .A1(b[0]), .A2(n505), .ZN(\intadd_8/A[0] ) );
  AOI22_X1 U835 ( .A1(b[6]), .A2(n633), .B1(n1), .B2(n764), .ZN(n506) );
  OAI221_X1 U836 ( .B1(b[5]), .B2(n631), .C1(n741), .C2(n643), .A(n506), .ZN(
        \intadd_8/B[0] ) );
  OAI221_X1 U837 ( .B1(a[1]), .B2(b[8]), .C1(n1239), .C2(n654), .A(a[0]), .ZN(
        n507) );
  OAI21_X1 U838 ( .B1(b[7]), .B2(n508), .A(n507), .ZN(\intadd_8/CI ) );
  FA_X1 U839 ( .A(n511), .B(n510), .CI(n509), .CO(n207), .S(\intadd_8/B[1] )
         );
  NAND2_X1 U840 ( .A1(n530), .A2(n704), .ZN(n512) );
  OAI221_X1 U841 ( .B1(b[5]), .B2(n527), .C1(n741), .C2(n528), .A(n512), .ZN(
        \intadd_26/A[0] ) );
  AOI22_X1 U842 ( .A1(b[1]), .A2(n715), .B1(n714), .B2(n628), .ZN(n513) );
  AOI221_X1 U843 ( .B1(n729), .B2(b[0]), .C1(n717), .C2(n1238), .A(n513), .ZN(
        n516) );
  OAI21_X1 U844 ( .B1(n514), .B2(n1247), .A(\intadd_3/B[0] ), .ZN(n515) );
  NOR2_X1 U845 ( .A1(n516), .A2(n515), .ZN(n521) );
  AOI21_X1 U846 ( .B1(n516), .B2(n515), .A(n521), .ZN(\intadd_26/B[0] ) );
  AOI22_X1 U847 ( .A1(b[3]), .A2(n633), .B1(n1), .B2(n555), .ZN(n517) );
  OAI221_X1 U848 ( .B1(b[2]), .B2(n631), .C1(n606), .C2(n643), .A(n517), .ZN(
        \intadd_26/CI ) );
  XOR2_X1 U849 ( .A(n519), .B(n518), .Z(n541) );
  XNOR2_X1 U850 ( .A(n540), .B(n541), .ZN(n524) );
  AOI22_X1 U851 ( .A1(b[4]), .A2(n633), .B1(n1), .B2(n704), .ZN(n520) );
  OAI221_X1 U852 ( .B1(b[3]), .B2(n631), .C1(n555), .C2(n643), .A(n520), .ZN(
        n522) );
  NOR2_X1 U853 ( .A1(n521), .A2(n522), .ZN(n539) );
  NOR2_X1 U854 ( .A1(n539), .A2(n537), .ZN(n523) );
  XNOR2_X1 U855 ( .A(n524), .B(n523), .ZN(\intadd_26/A[1] ) );
  AOI22_X1 U856 ( .A1(b[1]), .A2(n643), .B1(n631), .B2(n628), .ZN(n525) );
  AOI221_X1 U857 ( .B1(n633), .B2(b[2]), .C1(n1), .C2(n606), .A(n525), .ZN(
        n533) );
  NAND2_X1 U858 ( .A1(b[0]), .A2(n526), .ZN(n532) );
  AOI22_X1 U859 ( .A1(b[4]), .A2(n528), .B1(n527), .B2(n704), .ZN(n529) );
  AOI21_X1 U860 ( .B1(n530), .B2(n555), .A(n529), .ZN(n531) );
  FA_X1 U861 ( .A(n533), .B(n532), .CI(n531), .CO(n1047), .S(n1279) );
  OAI221_X1 U862 ( .B1(n534), .B2(n1274), .C1(n534), .C2(n1275), .A(n1277), 
        .ZN(n535) );
  NAND2_X1 U863 ( .A1(n1276), .A2(n535), .ZN(n1042) );
  INV_X1 U864 ( .A(\intadd_26/SUM[0] ), .ZN(n1046) );
  NOR3_X1 U865 ( .A1(n1274), .A2(n1275), .A3(n1277), .ZN(n1043) );
  OAI211_X1 U866 ( .C1(n1043), .C2(n1276), .A(n1045), .B(n535), .ZN(n536) );
  AOI22_X1 U867 ( .A1(n1047), .A2(n1042), .B1(n1046), .B2(n536), .ZN(
        \intadd_26/B[1] ) );
  NOR3_X1 U868 ( .A1(n541), .A2(n537), .A3(n540), .ZN(n538) );
  AOI211_X1 U869 ( .C1(n541), .C2(n540), .A(n539), .B(n538), .ZN(
        \intadd_26/B[2] ) );
  FA_X1 U870 ( .A(\intadd_28/SUM[0] ), .B(n543), .CI(n542), .CO(
        \intadd_8/B[4] ), .S(n218) );
  FA_X1 U871 ( .A(\intadd_21/n1 ), .B(\intadd_9/SUM[3] ), .CI(
        \intadd_10/SUM[2] ), .CO(\intadd_11/A[1] ), .S(\intadd_11/B[0] ) );
  AOI22_X1 U872 ( .A1(b[23]), .A2(n723), .B1(n773), .B2(n1151), .ZN(n544) );
  AOI221_X1 U873 ( .B1(n776), .B2(b[22]), .C1(n725), .C2(n1140), .A(n544), 
        .ZN(\intadd_25/A[0] ) );
  AOI22_X1 U874 ( .A1(b[9]), .A2(n1103), .B1(n1104), .B2(n689), .ZN(n545) );
  AOI221_X1 U875 ( .B1(n1101), .B2(b[8]), .C1(n1100), .C2(n654), .A(n545), 
        .ZN(\intadd_25/B[0] ) );
  AOI22_X1 U876 ( .A1(b[10]), .A2(n884), .B1(n885), .B2(n649), .ZN(n546) );
  AOI221_X1 U877 ( .B1(n882), .B2(b[11]), .C1(n881), .C2(n754), .A(n546), .ZN(
        \intadd_25/CI ) );
  AOI22_X1 U878 ( .A1(b[14]), .A2(n691), .B1(n690), .B2(n554), .ZN(n547) );
  AOI221_X1 U879 ( .B1(n694), .B2(b[15]), .C1(n693), .C2(n687), .A(n547), .ZN(
        \intadd_3/A[0] ) );
  AOI22_X1 U880 ( .A1(b[6]), .A2(n1150), .B1(n1108), .B2(n764), .ZN(n548) );
  AOI221_X1 U881 ( .B1(n1147), .B2(n712), .C1(n1139), .C2(b[7]), .A(n548), 
        .ZN(\intadd_3/CI ) );
  NOR2_X1 U882 ( .A1(n1105), .A2(n704), .ZN(n735) );
  AOI22_X1 U883 ( .A1(b[16]), .A2(n816), .B1(n815), .B2(n575), .ZN(n549) );
  OAI221_X1 U884 ( .B1(b[17]), .B2(n812), .C1(n824), .C2(n813), .A(n549), .ZN(
        n743) );
  AOI21_X1 U885 ( .B1(n704), .B2(n741), .A(n1105), .ZN(n739) );
  AOI22_X1 U886 ( .A1(b[5]), .A2(n735), .B1(n743), .B2(n739), .ZN(
        \intadd_3/A[1] ) );
  AOI22_X1 U887 ( .A1(b[15]), .A2(n691), .B1(n690), .B2(n687), .ZN(n550) );
  AOI221_X1 U888 ( .B1(n694), .B2(b[16]), .C1(n693), .C2(n575), .A(n550), .ZN(
        \intadd_3/B[1] ) );
  AOI22_X1 U889 ( .A1(b[16]), .A2(n813), .B1(n812), .B2(n575), .ZN(n551) );
  AOI221_X1 U890 ( .B1(n816), .B2(b[15]), .C1(n815), .C2(n687), .A(n551), .ZN(
        n560) );
  AOI22_X1 U891 ( .A1(b[13]), .A2(n691), .B1(n690), .B2(n637), .ZN(n552) );
  AOI221_X1 U892 ( .B1(n694), .B2(b[14]), .C1(n693), .C2(n554), .A(n552), .ZN(
        n559) );
  NAND2_X1 U893 ( .A1(n560), .A2(n559), .ZN(n569) );
  AOI22_X1 U894 ( .A1(b[15]), .A2(n813), .B1(n812), .B2(n687), .ZN(n553) );
  AOI221_X1 U895 ( .B1(n816), .B2(b[14]), .C1(n815), .C2(n554), .A(n553), .ZN(
        n710) );
  NOR2_X1 U896 ( .A1(n1105), .A2(n555), .ZN(n703) );
  OAI21_X1 U897 ( .B1(a[23]), .B2(b[4]), .A(n740), .ZN(n577) );
  OAI22_X1 U898 ( .A1(b[5]), .A2(n604), .B1(n605), .B2(n577), .ZN(n556) );
  AOI211_X1 U899 ( .C1(b[5]), .C2(n1139), .A(n703), .B(n556), .ZN(n558) );
  NAND2_X1 U900 ( .A1(n703), .A2(n556), .ZN(n557) );
  OAI21_X1 U901 ( .B1(n710), .B2(n558), .A(n557), .ZN(n573) );
  NOR2_X1 U902 ( .A1(n560), .A2(n559), .ZN(n571) );
  AOI21_X1 U903 ( .B1(n569), .B2(n573), .A(n571), .ZN(\intadd_17/B[2] ) );
  AOI22_X1 U904 ( .A1(b[11]), .A2(n826), .B1(n825), .B2(n754), .ZN(n561) );
  AOI221_X1 U905 ( .B1(n846), .B2(b[10]), .C1(n828), .C2(n649), .A(n561), .ZN(
        \intadd_17/A[0] ) );
  AOI22_X1 U906 ( .A1(b[8]), .A2(n884), .B1(n885), .B2(n654), .ZN(n562) );
  AOI221_X1 U907 ( .B1(n882), .B2(b[9]), .C1(n881), .C2(n689), .A(n562), .ZN(
        \intadd_17/B[0] ) );
  AOI22_X1 U908 ( .A1(b[19]), .A2(n780), .B1(n720), .B2(n1106), .ZN(n563) );
  AOI221_X1 U909 ( .B1(n771), .B2(b[18]), .C1(n722), .C2(n1114), .A(n563), 
        .ZN(\intadd_17/CI ) );
  AOI22_X1 U910 ( .A1(b[13]), .A2(n694), .B1(n693), .B2(n637), .ZN(n564) );
  OAI221_X1 U911 ( .B1(b[12]), .B2(n690), .C1(n650), .C2(n691), .A(n564), .ZN(
        n862) );
  NOR3_X1 U912 ( .A1(n1239), .A2(n565), .A3(a[2]), .ZN(n664) );
  INV_X1 U913 ( .A(n664), .ZN(n659) );
  NOR2_X1 U914 ( .A1(a[1]), .A2(a[3]), .ZN(n585) );
  AOI21_X1 U915 ( .B1(n862), .B2(n659), .A(n585), .ZN(\intadd_17/B[1] ) );
  AOI22_X1 U916 ( .A1(b[9]), .A2(n884), .B1(n885), .B2(n689), .ZN(n566) );
  AOI221_X1 U917 ( .B1(n882), .B2(b[10]), .C1(n881), .C2(n649), .A(n566), .ZN(
        \intadd_4/A[0] ) );
  AOI22_X1 U918 ( .A1(b[8]), .A2(n1103), .B1(n1104), .B2(n654), .ZN(n567) );
  AOI221_X1 U919 ( .B1(n1101), .B2(b[7]), .C1(n1100), .C2(n712), .A(n567), 
        .ZN(\intadd_4/B[0] ) );
  AOI22_X1 U920 ( .A1(b[12]), .A2(n826), .B1(n825), .B2(n650), .ZN(n568) );
  AOI221_X1 U921 ( .B1(n846), .B2(b[11]), .C1(n828), .C2(n754), .A(n568), .ZN(
        \intadd_4/CI ) );
  NOR2_X1 U922 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U923 ( .A(n573), .B(n572), .ZN(\intadd_15/A[2] ) );
  AOI22_X1 U924 ( .A1(b[17]), .A2(n791), .B1(n790), .B2(n824), .ZN(n574) );
  AOI221_X1 U925 ( .B1(n819), .B2(b[16]), .C1(n793), .C2(n575), .A(n574), .ZN(
        \intadd_15/A[1] ) );
  OAI22_X1 U926 ( .A1(b[3]), .A2(n1108), .B1(n577), .B2(n576), .ZN(n578) );
  AOI21_X1 U927 ( .B1(b[3]), .B2(n1138), .A(n578), .ZN(\intadd_15/A[0] ) );
  AOI22_X1 U928 ( .A1(b[5]), .A2(n624), .B1(n623), .B2(n741), .ZN(n579) );
  AOI221_X1 U929 ( .B1(n626), .B2(b[6]), .C1(n1096), .C2(n764), .A(n579), .ZN(
        \intadd_15/B[0] ) );
  AOI221_X1 U930 ( .B1(\intadd_3/B[0] ), .B2(n1140), .C1(n726), .C2(b[22]), 
        .A(n717), .ZN(n582) );
  AOI22_X1 U931 ( .A1(n582), .A2(n581), .B1(n580), .B2(n878), .ZN(n583) );
  OAI221_X1 U932 ( .B1(n584), .B2(a[5]), .C1(n584), .C2(n878), .A(n583), .ZN(
        \intadd_15/CI ) );
  NOR2_X1 U933 ( .A1(n1105), .A2(n606), .ZN(n668) );
  OAI211_X1 U934 ( .C1(n662), .C2(n1151), .A(n659), .B(n666), .ZN(n586) );
  OAI211_X1 U935 ( .C1(n661), .C2(n1151), .A(n663), .B(n586), .ZN(
        \intadd_15/B[1] ) );
  AOI22_X1 U936 ( .A1(b[10]), .A2(n1103), .B1(n1104), .B2(n649), .ZN(n587) );
  AOI221_X1 U937 ( .B1(n1101), .B2(b[9]), .C1(n1100), .C2(n689), .A(n587), 
        .ZN(\intadd_1/A[0] ) );
  AOI22_X1 U938 ( .A1(b[20]), .A2(n791), .B1(n790), .B2(n1098), .ZN(n588) );
  AOI221_X1 U939 ( .B1(n819), .B2(b[19]), .C1(n793), .C2(n1106), .A(n588), 
        .ZN(\intadd_1/B[0] ) );
  AOI22_X1 U940 ( .A1(b[7]), .A2(n1150), .B1(n1108), .B2(n712), .ZN(n589) );
  AOI221_X1 U941 ( .B1(n1147), .B2(n654), .C1(n1139), .C2(b[8]), .A(n589), 
        .ZN(\intadd_1/CI ) );
  AOI21_X1 U942 ( .B1(n712), .B2(n764), .A(n1105), .ZN(n766) );
  OAI21_X1 U943 ( .B1(n764), .B2(n712), .A(n766), .ZN(n591) );
  AOI22_X1 U944 ( .A1(b[17]), .A2(n694), .B1(n693), .B2(n824), .ZN(n590) );
  OAI221_X1 U945 ( .B1(b[16]), .B2(n690), .C1(n575), .C2(n691), .A(n590), .ZN(
        n765) );
  XOR2_X1 U946 ( .A(n591), .B(n765), .Z(\intadd_1/A[1] ) );
  AOI22_X1 U947 ( .A1(b[11]), .A2(n884), .B1(n885), .B2(n754), .ZN(n592) );
  AOI221_X1 U948 ( .B1(n882), .B2(b[12]), .C1(n881), .C2(n650), .A(n592), .ZN(
        n597) );
  AOI22_X1 U949 ( .A1(b[18]), .A2(n813), .B1(n812), .B2(n1114), .ZN(n593) );
  AOI221_X1 U950 ( .B1(n816), .B2(b[17]), .C1(n815), .C2(n824), .A(n593), .ZN(
        n596) );
  AOI22_X1 U951 ( .A1(b[14]), .A2(n826), .B1(n825), .B2(n554), .ZN(n594) );
  AOI221_X1 U952 ( .B1(n846), .B2(b[13]), .C1(n828), .C2(n637), .A(n594), .ZN(
        n595) );
  FA_X1 U953 ( .A(n597), .B(n596), .CI(n595), .CO(\intadd_1/B[1] ), .S(
        \intadd_4/B[2] ) );
  AOI22_X1 U954 ( .A1(b[19]), .A2(n813), .B1(n812), .B2(n1106), .ZN(n598) );
  AOI221_X1 U955 ( .B1(n816), .B2(b[18]), .C1(n815), .C2(n1114), .A(n598), 
        .ZN(\intadd_2/A[0] ) );
  AOI22_X1 U956 ( .A1(b[12]), .A2(n884), .B1(n885), .B2(n650), .ZN(n599) );
  AOI221_X1 U957 ( .B1(n882), .B2(b[13]), .C1(n881), .C2(n637), .A(n599), .ZN(
        \intadd_2/B[0] ) );
  AOI22_X1 U958 ( .A1(b[11]), .A2(n1103), .B1(n1104), .B2(n754), .ZN(n600) );
  AOI221_X1 U959 ( .B1(n1101), .B2(b[10]), .C1(n1100), .C2(n649), .A(n600), 
        .ZN(\intadd_2/CI ) );
  AOI22_X1 U960 ( .A1(b[21]), .A2(n780), .B1(n720), .B2(n878), .ZN(n601) );
  AOI221_X1 U961 ( .B1(n771), .B2(b[20]), .C1(n722), .C2(n1098), .A(n601), 
        .ZN(n738) );
  AOI22_X1 U962 ( .A1(b[19]), .A2(n791), .B1(n790), .B2(n1106), .ZN(n602) );
  AOI221_X1 U963 ( .B1(n819), .B2(b[18]), .C1(n793), .C2(n1114), .A(n602), 
        .ZN(n737) );
  AOI22_X1 U964 ( .A1(b[13]), .A2(n826), .B1(n825), .B2(n637), .ZN(n603) );
  AOI221_X1 U965 ( .B1(n846), .B2(b[12]), .C1(n828), .C2(n650), .A(n603), .ZN(
        n736) );
  NOR2_X1 U966 ( .A1(b[3]), .A2(n604), .ZN(n708) );
  AOI211_X1 U967 ( .C1(n1105), .C2(n606), .A(n668), .B(n605), .ZN(n607) );
  AOI211_X1 U968 ( .C1(n1139), .C2(b[3]), .A(n708), .B(n607), .ZN(
        \intadd_5/A[0] ) );
  AOI22_X1 U969 ( .A1(b[5]), .A2(n1103), .B1(n1104), .B2(n741), .ZN(n608) );
  AOI221_X1 U970 ( .B1(n1101), .B2(b[4]), .C1(n1100), .C2(n704), .A(n608), 
        .ZN(\intadd_5/B[0] ) );
  AOI22_X1 U971 ( .A1(b[21]), .A2(n715), .B1(n714), .B2(n878), .ZN(n609) );
  AOI221_X1 U972 ( .B1(n729), .B2(b[20]), .C1(n717), .C2(n1098), .A(n609), 
        .ZN(\intadd_5/CI ) );
  FA_X1 U973 ( .A(n612), .B(n611), .CI(n610), .CO(n617), .S(n394) );
  OAI21_X1 U974 ( .B1(b[1]), .B2(n1105), .A(n1108), .ZN(n613) );
  NAND3_X1 U975 ( .A1(n1247), .A2(n1164), .A3(n613), .ZN(n616) );
  AOI22_X1 U976 ( .A1(b[14]), .A2(n791), .B1(n790), .B2(n554), .ZN(n614) );
  AOI221_X1 U977 ( .B1(n819), .B2(b[13]), .C1(n793), .C2(n637), .A(n614), .ZN(
        n615) );
  FA_X1 U978 ( .A(n617), .B(n616), .CI(n615), .CO(\intadd_16/B[2] ), .S(
        \intadd_24/B[2] ) );
  AOI22_X1 U979 ( .A1(b[14]), .A2(n813), .B1(n812), .B2(n554), .ZN(n618) );
  AOI221_X1 U980 ( .B1(n816), .B2(b[13]), .C1(n815), .C2(n637), .A(n618), .ZN(
        \intadd_5/A[1] ) );
  NOR2_X1 U981 ( .A1(n1105), .A2(n628), .ZN(n645) );
  INV_X1 U982 ( .A(n645), .ZN(n619) );
  AOI221_X1 U983 ( .B1(n1140), .B2(n619), .C1(n662), .C2(n619), .A(n1239), 
        .ZN(n622) );
  NOR2_X1 U984 ( .A1(b[22]), .A2(n631), .ZN(n620) );
  AOI221_X1 U985 ( .B1(n633), .B2(b[23]), .C1(n1), .C2(n1163), .A(n620), .ZN(
        n642) );
  INV_X1 U986 ( .A(n642), .ZN(n621) );
  OAI22_X1 U987 ( .A1(a[1]), .A2(n645), .B1(n622), .B2(n621), .ZN(
        \intadd_5/B[1] ) );
  OAI21_X1 U988 ( .B1(a[0]), .B2(n1151), .A(a[1]), .ZN(n635) );
  AOI22_X1 U989 ( .A1(b[3]), .A2(n624), .B1(n623), .B2(n555), .ZN(n625) );
  AOI221_X1 U990 ( .B1(n626), .B2(b[4]), .C1(n1096), .C2(n704), .A(n625), .ZN(
        n634) );
  AOI22_X1 U991 ( .A1(b[5]), .A2(n884), .B1(n885), .B2(n741), .ZN(n627) );
  AOI221_X1 U992 ( .B1(n882), .B2(b[6]), .C1(n881), .C2(n764), .A(n627), .ZN(
        n675) );
  AOI21_X1 U993 ( .B1(n1105), .B2(n606), .A(n668), .ZN(n630) );
  AOI22_X1 U994 ( .A1(b[1]), .A2(n1150), .B1(n1108), .B2(n628), .ZN(n629) );
  AOI21_X1 U995 ( .B1(n701), .B2(n630), .A(n629), .ZN(n674) );
  AOI22_X1 U996 ( .A1(b[21]), .A2(n643), .B1(n631), .B2(n878), .ZN(n632) );
  AOI221_X1 U997 ( .B1(n633), .B2(b[22]), .C1(n1), .C2(n1140), .A(n632), .ZN(
        n673) );
  FA_X1 U998 ( .A(n636), .B(n635), .CI(n634), .CO(n640), .S(\intadd_16/B[1] )
         );
  AOI22_X1 U999 ( .A1(b[13]), .A2(n813), .B1(n812), .B2(n637), .ZN(n638) );
  AOI221_X1 U1000 ( .B1(n816), .B2(b[12]), .C1(n815), .C2(n650), .A(n638), 
        .ZN(n639) );
  FA_X1 U1001 ( .A(n641), .B(n640), .CI(n639), .CO(\intadd_27/B[2] ), .S(
        \intadd_16/A[2] ) );
  OAI21_X1 U1002 ( .B1(n1140), .B2(n643), .A(n642), .ZN(n644) );
  XNOR2_X1 U1003 ( .A(a[1]), .B(n644), .ZN(n646) );
  XOR2_X1 U1004 ( .A(n646), .B(n645), .Z(\intadd_27/B[1] ) );
  AOI22_X1 U1005 ( .A1(b[16]), .A2(n780), .B1(n720), .B2(n575), .ZN(n647) );
  AOI221_X1 U1006 ( .B1(n771), .B2(b[15]), .C1(n722), .C2(n687), .A(n647), 
        .ZN(n672) );
  AOI22_X1 U1007 ( .A1(b[9]), .A2(n691), .B1(n690), .B2(n689), .ZN(n648) );
  AOI221_X1 U1008 ( .B1(n694), .B2(b[10]), .C1(n693), .C2(n649), .A(n648), 
        .ZN(n671) );
  AOI22_X1 U1009 ( .A1(b[12]), .A2(n813), .B1(n812), .B2(n650), .ZN(n651) );
  AOI221_X1 U1010 ( .B1(n816), .B2(b[11]), .C1(n815), .C2(n754), .A(n651), 
        .ZN(n670) );
  AOI22_X1 U1011 ( .A1(b[10]), .A2(n691), .B1(n690), .B2(n649), .ZN(n652) );
  AOI221_X1 U1012 ( .B1(n694), .B2(b[11]), .C1(n693), .C2(n754), .A(n652), 
        .ZN(n683) );
  AOI22_X1 U1013 ( .A1(b[9]), .A2(n826), .B1(n825), .B2(n689), .ZN(n653) );
  AOI221_X1 U1014 ( .B1(n846), .B2(b[8]), .C1(n828), .C2(n654), .A(n653), .ZN(
        n682) );
  AOI22_X1 U1015 ( .A1(b[15]), .A2(n791), .B1(n790), .B2(n687), .ZN(n655) );
  AOI221_X1 U1016 ( .B1(n819), .B2(b[14]), .C1(n793), .C2(n554), .A(n655), 
        .ZN(n681) );
  AOI22_X1 U1017 ( .A1(b[17]), .A2(n780), .B1(n720), .B2(n824), .ZN(n656) );
  AOI221_X1 U1018 ( .B1(n771), .B2(b[16]), .C1(n722), .C2(n575), .A(n656), 
        .ZN(n680) );
  AOI22_X1 U1019 ( .A1(b[19]), .A2(n723), .B1(n773), .B2(n1106), .ZN(n657) );
  AOI221_X1 U1020 ( .B1(n776), .B2(b[18]), .C1(n725), .C2(n1114), .A(n657), 
        .ZN(n679) );
  AOI22_X1 U1021 ( .A1(b[6]), .A2(n884), .B1(n885), .B2(n764), .ZN(n658) );
  AOI221_X1 U1022 ( .B1(n882), .B2(b[7]), .C1(n881), .C2(n712), .A(n658), .ZN(
        n678) );
  NAND2_X1 U1023 ( .A1(n662), .A2(n661), .ZN(n660) );
  NAND2_X1 U1024 ( .A1(n663), .A2(n659), .ZN(n863) );
  AOI21_X1 U1025 ( .B1(b[23]), .B2(n660), .A(n863), .ZN(n669) );
  AOI22_X1 U1026 ( .A1(n1151), .A2(n663), .B1(n662), .B2(n661), .ZN(n665) );
  OR3_X1 U1027 ( .A1(n666), .A2(n665), .A3(n664), .ZN(n667) );
  OAI21_X1 U1028 ( .B1(n669), .B2(n668), .A(n667), .ZN(n868) );
  FA_X1 U1029 ( .A(n672), .B(n671), .CI(n670), .CO(\intadd_27/A[1] ), .S(n677)
         );
  FA_X1 U1030 ( .A(n675), .B(n674), .CI(n673), .CO(n641), .S(n676) );
  FA_X1 U1031 ( .A(\intadd_27/SUM[0] ), .B(n677), .CI(n676), .CO(n685), .S(
        \intadd_6/A[2] ) );
  FA_X1 U1032 ( .A(n680), .B(n679), .CI(n678), .CO(n869), .S(n867) );
  FA_X1 U1033 ( .A(n683), .B(n682), .CI(n681), .CO(n870), .S(n866) );
  FA_X1 U1034 ( .A(\intadd_27/SUM[1] ), .B(n685), .CI(n684), .CO(
        \intadd_16/B[3] ), .S(\intadd_7/A[4] ) );
  AOI22_X1 U1035 ( .A1(b[16]), .A2(n791), .B1(n790), .B2(n575), .ZN(n686) );
  AOI221_X1 U1036 ( .B1(n819), .B2(b[15]), .C1(n793), .C2(n687), .A(n686), 
        .ZN(n855) );
  AOI22_X1 U1037 ( .A1(b[10]), .A2(n826), .B1(n825), .B2(n649), .ZN(n688) );
  AOI221_X1 U1038 ( .B1(n846), .B2(b[9]), .C1(n828), .C2(n689), .A(n688), .ZN(
        n854) );
  AOI22_X1 U1039 ( .A1(b[11]), .A2(n691), .B1(n690), .B2(n754), .ZN(n692) );
  AOI221_X1 U1040 ( .B1(n694), .B2(b[12]), .C1(n693), .C2(n650), .A(n692), 
        .ZN(n853) );
  NAND3_X1 U1041 ( .A1(a[7]), .A2(b[17]), .A3(n767), .ZN(n696) );
  AOI221_X1 U1042 ( .B1(a[9]), .B2(n1114), .C1(n767), .C2(b[18]), .A(n771), 
        .ZN(n695) );
  AOI21_X1 U1043 ( .B1(n768), .B2(n696), .A(n695), .ZN(n697) );
  AOI21_X1 U1044 ( .B1(n722), .B2(n824), .A(n697), .ZN(n858) );
  AOI22_X1 U1045 ( .A1(b[20]), .A2(n723), .B1(n773), .B2(n1098), .ZN(n698) );
  AOI221_X1 U1046 ( .B1(n776), .B2(b[19]), .C1(n725), .C2(n1106), .A(n698), 
        .ZN(n857) );
  AOI22_X1 U1047 ( .A1(b[7]), .A2(n884), .B1(n885), .B2(n712), .ZN(n699) );
  AOI221_X1 U1048 ( .B1(n882), .B2(b[8]), .C1(n881), .C2(n654), .A(n699), .ZN(
        n856) );
  NOR2_X1 U1049 ( .A1(a[21]), .A2(a[22]), .ZN(n700) );
  AOI22_X1 U1050 ( .A1(n701), .A2(n741), .B1(n700), .B2(n704), .ZN(n702) );
  NOR2_X1 U1051 ( .A1(n702), .A2(n555), .ZN(n706) );
  AOI21_X1 U1052 ( .B1(n1141), .B2(n704), .A(n703), .ZN(n705) );
  OAI22_X1 U1053 ( .A1(n706), .A2(n705), .B1(n704), .B2(n1150), .ZN(n707) );
  AOI221_X1 U1054 ( .B1(n1139), .B2(b[5]), .C1(n708), .C2(n741), .A(n707), 
        .ZN(n709) );
  XNOR2_X1 U1055 ( .A(n710), .B(n709), .ZN(n850) );
  AOI22_X1 U1056 ( .A1(b[21]), .A2(n723), .B1(n773), .B2(n878), .ZN(n711) );
  AOI221_X1 U1057 ( .B1(n776), .B2(b[20]), .C1(n725), .C2(n1098), .A(n711), 
        .ZN(n861) );
  AOI22_X1 U1058 ( .A1(b[7]), .A2(n1103), .B1(n1104), .B2(n712), .ZN(n713) );
  AOI221_X1 U1059 ( .B1(n1101), .B2(b[6]), .C1(n1100), .C2(n764), .A(n713), 
        .ZN(n860) );
  AOI22_X1 U1060 ( .A1(b[23]), .A2(n715), .B1(n714), .B2(n1151), .ZN(n716) );
  AOI221_X1 U1061 ( .B1(n729), .B2(b[22]), .C1(n717), .C2(n1140), .A(n716), 
        .ZN(n859) );
  AOI22_X1 U1062 ( .A1(b[5]), .A2(n1150), .B1(n1108), .B2(n741), .ZN(n718) );
  AOI221_X1 U1063 ( .B1(n1147), .B2(n764), .C1(n1139), .C2(b[6]), .A(n718), 
        .ZN(n732) );
  AOI22_X1 U1064 ( .A1(b[18]), .A2(n791), .B1(n790), .B2(n1114), .ZN(n719) );
  AOI221_X1 U1065 ( .B1(n819), .B2(b[17]), .C1(n793), .C2(n824), .A(n719), 
        .ZN(n731) );
  AOI22_X1 U1066 ( .A1(b[20]), .A2(n780), .B1(n720), .B2(n1098), .ZN(n721) );
  AOI221_X1 U1067 ( .B1(n771), .B2(b[19]), .C1(n722), .C2(n1106), .A(n721), 
        .ZN(n730) );
  AOI22_X1 U1068 ( .A1(b[22]), .A2(n723), .B1(n773), .B2(n1140), .ZN(n724) );
  AOI221_X1 U1069 ( .B1(n776), .B2(b[21]), .C1(n725), .C2(n878), .A(n724), 
        .ZN(n734) );
  NOR2_X1 U1070 ( .A1(a[3]), .A2(n726), .ZN(n728) );
  AOI221_X1 U1071 ( .B1(n729), .B2(b[23]), .C1(n728), .C2(n1163), .A(n727), 
        .ZN(n733) );
  FA_X1 U1072 ( .A(n732), .B(n731), .CI(n730), .CO(\intadd_4/B[1] ), .S(n872)
         );
  FA_X1 U1073 ( .A(n735), .B(n734), .CI(n733), .CO(\intadd_4/A[1] ), .S(n871)
         );
  FA_X1 U1074 ( .A(n738), .B(n737), .CI(n736), .CO(\intadd_25/B[1] ), .S(n849)
         );
  OAI21_X1 U1075 ( .B1(n741), .B2(n740), .A(n739), .ZN(n742) );
  XOR2_X1 U1076 ( .A(n743), .B(n742), .Z(n848) );
  FA_X1 U1077 ( .A(\intadd_4/SUM[1] ), .B(n745), .CI(n744), .CO(
        \intadd_17/B[3] ), .S(\intadd_5/B[4] ) );
  FA_X1 U1078 ( .A(n748), .B(n747), .CI(n746), .CO(n146), .S(n758) );
  FA_X1 U1079 ( .A(n751), .B(n750), .CI(n749), .CO(n798), .S(n757) );
  AOI22_X1 U1080 ( .A1(b[13]), .A2(n884), .B1(n885), .B2(n637), .ZN(n752) );
  AOI221_X1 U1081 ( .B1(n882), .B2(b[14]), .C1(n881), .C2(n554), .A(n752), 
        .ZN(n835) );
  AOI22_X1 U1082 ( .A1(b[12]), .A2(n1103), .B1(n1104), .B2(n650), .ZN(n753) );
  AOI221_X1 U1083 ( .B1(n1101), .B2(b[11]), .C1(n1100), .C2(n754), .A(n753), 
        .ZN(n834) );
  AOI22_X1 U1084 ( .A1(b[16]), .A2(n826), .B1(n825), .B2(n575), .ZN(n755) );
  AOI221_X1 U1085 ( .B1(n846), .B2(b[15]), .C1(n828), .C2(n687), .A(n755), 
        .ZN(n833) );
  FA_X1 U1086 ( .A(n758), .B(n757), .CI(n756), .CO(\intadd_1/A[3] ), .S(
        \intadd_3/A[3] ) );
  AOI22_X1 U1087 ( .A1(b[8]), .A2(n1150), .B1(n1108), .B2(n654), .ZN(n759) );
  AOI221_X1 U1088 ( .B1(n1147), .B2(n689), .C1(n1139), .C2(b[9]), .A(n759), 
        .ZN(n763) );
  AOI22_X1 U1089 ( .A1(b[15]), .A2(n826), .B1(n825), .B2(n687), .ZN(n760) );
  AOI221_X1 U1090 ( .B1(n846), .B2(b[14]), .C1(n828), .C2(n554), .A(n760), 
        .ZN(n762) );
  FA_X1 U1091 ( .A(n763), .B(n762), .CI(n761), .CO(\intadd_2/A[1] ), .S(
        \intadd_3/A[2] ) );
  NOR2_X1 U1092 ( .A1(n1105), .A2(n764), .ZN(n777) );
  AOI22_X1 U1093 ( .A1(b[7]), .A2(n777), .B1(n766), .B2(n765), .ZN(
        \intadd_2/B[1] ) );
  AOI22_X1 U1094 ( .A1(b[22]), .A2(n767), .B1(a[9]), .B2(n1140), .ZN(n781) );
  OAI22_X1 U1095 ( .A1(b[21]), .A2(n769), .B1(n768), .B2(n781), .ZN(n770) );
  AOI21_X1 U1096 ( .B1(n771), .B2(b[21]), .A(n770), .ZN(n779) );
  NOR2_X1 U1097 ( .A1(a[6]), .A2(n772), .ZN(n775) );
  AOI221_X1 U1098 ( .B1(n776), .B2(b[23]), .C1(n775), .C2(n1163), .A(n774), 
        .ZN(n778) );
  FA_X1 U1099 ( .A(n779), .B(n778), .CI(n777), .CO(n788), .S(\intadd_25/A[1] )
         );
  OAI22_X1 U1100 ( .A1(n782), .A2(n781), .B1(n1151), .B2(n780), .ZN(n783) );
  AOI21_X1 U1101 ( .B1(n784), .B2(n1151), .A(n783), .ZN(n787) );
  AOI22_X1 U1102 ( .A1(b[21]), .A2(n791), .B1(n790), .B2(n878), .ZN(n785) );
  AOI221_X1 U1103 ( .B1(n819), .B2(b[20]), .C1(n793), .C2(n1098), .A(n785), 
        .ZN(n786) );
  FA_X1 U1104 ( .A(n788), .B(n787), .CI(n786), .CO(\intadd_1/B[2] ), .S(
        \intadd_25/B[2] ) );
  AOI22_X1 U1105 ( .A1(b[14]), .A2(n884), .B1(n885), .B2(n554), .ZN(n789) );
  AOI221_X1 U1106 ( .B1(n882), .B2(b[15]), .C1(n881), .C2(n687), .A(n789), 
        .ZN(\intadd_13/A[0] ) );
  AOI22_X1 U1107 ( .A1(b[23]), .A2(n791), .B1(n790), .B2(n1151), .ZN(n792) );
  AOI221_X1 U1108 ( .B1(n819), .B2(b[22]), .C1(n793), .C2(n1140), .A(n792), 
        .ZN(\intadd_13/B[0] ) );
  AOI22_X1 U1109 ( .A1(b[13]), .A2(n1103), .B1(n1104), .B2(n637), .ZN(n794) );
  AOI221_X1 U1110 ( .B1(n1101), .B2(b[12]), .C1(n1100), .C2(n650), .A(n794), 
        .ZN(\intadd_13/CI ) );
  NAND2_X1 U1111 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U1112 ( .A(n798), .B(n797), .ZN(\intadd_2/B[2] ) );
  FA_X1 U1113 ( .A(n800), .B(\intadd_35/SUM[0] ), .CI(n799), .CO(n889), .S(
        \intadd_13/B[3] ) );
  FA_X1 U1114 ( .A(n803), .B(n802), .CI(n801), .CO(n811), .S(n135) );
  FA_X1 U1115 ( .A(n806), .B(n805), .CI(n804), .CO(n800), .S(n810) );
  FA_X1 U1116 ( .A(n818), .B(n808), .CI(n807), .CO(n282), .S(n809) );
  FA_X1 U1117 ( .A(n811), .B(n810), .CI(n809), .CO(\intadd_14/A[2] ), .S(
        \intadd_13/A[2] ) );
  AOI22_X1 U1118 ( .A1(b[22]), .A2(n813), .B1(n812), .B2(n1140), .ZN(n814) );
  AOI221_X1 U1119 ( .B1(n816), .B2(b[21]), .C1(n815), .C2(n878), .A(n814), 
        .ZN(n822) );
  NOR2_X1 U1120 ( .A1(n1105), .A2(n649), .ZN(n821) );
  AOI221_X1 U1121 ( .B1(n819), .B2(b[23]), .C1(n818), .C2(n1163), .A(n817), 
        .ZN(n820) );
  FA_X1 U1122 ( .A(n822), .B(n821), .CI(n820), .CO(\intadd_14/A[1] ), .S(
        \intadd_13/A[1] ) );
  AOI22_X1 U1123 ( .A1(b[10]), .A2(n1150), .B1(n1108), .B2(n649), .ZN(n823) );
  AOI221_X1 U1124 ( .B1(n1139), .B2(b[11]), .C1(n1147), .C2(n754), .A(n823), 
        .ZN(n832) );
  AOI22_X1 U1125 ( .A1(b[17]), .A2(n826), .B1(n825), .B2(n824), .ZN(n827) );
  AOI221_X1 U1126 ( .B1(n846), .B2(b[16]), .C1(n828), .C2(n575), .A(n827), 
        .ZN(n831) );
  FA_X1 U1127 ( .A(n832), .B(n831), .CI(n830), .CO(\intadd_13/B[1] ), .S(
        \intadd_2/A[2] ) );
  FA_X1 U1128 ( .A(n835), .B(n834), .CI(n833), .CO(n840), .S(n756) );
  OAI21_X1 U1129 ( .B1(n654), .B2(n689), .A(n836), .ZN(n837) );
  XOR2_X1 U1130 ( .A(n838), .B(n837), .Z(n839) );
  FA_X1 U1131 ( .A(n840), .B(\intadd_13/SUM[0] ), .CI(n839), .CO(
        \intadd_2/B[3] ), .S(\intadd_1/B[3] ) );
  AOI22_X1 U1132 ( .A1(b[22]), .A2(n1103), .B1(n1104), .B2(n1140), .ZN(n841)
         );
  AOI221_X1 U1133 ( .B1(n1101), .B2(b[21]), .C1(n1100), .C2(n878), .A(n841), 
        .ZN(\intadd_12/A[0] ) );
  NOR2_X1 U1134 ( .A1(n1114), .A2(n1105), .ZN(\intadd_12/B[0] ) );
  INV_X1 U1135 ( .A(n884), .ZN(n844) );
  NOR2_X1 U1136 ( .A1(a[17]), .A2(n842), .ZN(n843) );
  AOI221_X1 U1137 ( .B1(n844), .B2(b[23]), .C1(n843), .C2(n1163), .A(n881), 
        .ZN(\intadd_12/CI ) );
  AOI221_X1 U1138 ( .B1(n846), .B2(b[23]), .C1(n984), .C2(n1163), .A(n845), 
        .ZN(n877) );
  AOI22_X1 U1139 ( .A1(b[21]), .A2(n884), .B1(n885), .B2(n878), .ZN(n847) );
  AOI221_X1 U1140 ( .B1(n882), .B2(b[22]), .C1(n881), .C2(n1140), .A(n847), 
        .ZN(n876) );
  NOR2_X1 U1141 ( .A1(n1105), .A2(n575), .ZN(n875) );
  FA_X1 U1142 ( .A(n849), .B(n848), .CI(\intadd_25/SUM[0] ), .CO(n926), .S(
        n744) );
  FA_X1 U1143 ( .A(n852), .B(n851), .CI(n850), .CO(\intadd_15/B[2] ), .S(n930)
         );
  FA_X1 U1144 ( .A(n855), .B(n854), .CI(n853), .CO(n852), .S(n865) );
  FA_X1 U1145 ( .A(n858), .B(n857), .CI(n856), .CO(n851), .S(n864) );
  FA_X1 U1146 ( .A(n861), .B(n860), .CI(n859), .CO(\intadd_17/A[1] ), .S(n874)
         );
  XOR2_X1 U1147 ( .A(n863), .B(n862), .Z(n873) );
  FA_X1 U1148 ( .A(n865), .B(\intadd_15/SUM[0] ), .CI(n864), .CO(n929), .S(
        n933) );
  FA_X1 U1149 ( .A(n867), .B(n866), .CI(\intadd_5/SUM[0] ), .CO(n932), .S(n684) );
  FA_X1 U1150 ( .A(n870), .B(n869), .CI(n868), .CO(\intadd_5/B[2] ), .S(n931)
         );
  FA_X1 U1151 ( .A(n872), .B(n871), .CI(\intadd_4/SUM[0] ), .CO(n745), .S(n936) );
  FA_X1 U1152 ( .A(n874), .B(n873), .CI(\intadd_17/SUM[0] ), .CO(n935), .S(
        n928) );
  FA_X1 U1153 ( .A(n877), .B(n876), .CI(n875), .CO(n991), .S(\intadd_22/A[2] )
         );
  AOI22_X1 U1154 ( .A1(b[21]), .A2(n1103), .B1(n1104), .B2(n878), .ZN(n879) );
  AOI221_X1 U1155 ( .B1(n1101), .B2(b[20]), .C1(n1100), .C2(n1098), .A(n879), 
        .ZN(n983) );
  AOI22_X1 U1156 ( .A1(b[18]), .A2(n1150), .B1(n1108), .B2(n1114), .ZN(n880)
         );
  AOI221_X1 U1157 ( .B1(n1139), .B2(b[19]), .C1(n1147), .C2(n1106), .A(n880), 
        .ZN(n982) );
  AOI22_X1 U1158 ( .A1(b[23]), .A2(n882), .B1(n881), .B2(n1151), .ZN(n883) );
  OAI221_X1 U1159 ( .B1(b[22]), .B2(n885), .C1(n1140), .C2(n884), .A(n883), 
        .ZN(n986) );
  AOI21_X1 U1160 ( .B1(n575), .B2(n824), .A(n1105), .ZN(n985) );
  OAI21_X1 U1161 ( .B1(n575), .B2(n824), .A(n985), .ZN(n886) );
  XOR2_X1 U1162 ( .A(n986), .B(n886), .Z(n989) );
  INV_X1 U1163 ( .A(\intadd_23/SUM[1] ), .ZN(n893) );
  INV_X2 U1164 ( .A(\intadd_35/SUM[2] ), .ZN(n892) );
  AOI21_X1 U1165 ( .B1(n889), .B2(n888), .A(n887), .ZN(n891) );
  INV_X1 U1166 ( .A(n890), .ZN(n894) );
  NOR2_X1 U1167 ( .A1(n895), .A2(n894), .ZN(n1013) );
  INV_X1 U1168 ( .A(\intadd_14/n1 ), .ZN(n899) );
  FA_X1 U1169 ( .A(n893), .B(n892), .CI(n891), .CO(n890), .S(n900) );
  NOR2_X1 U1170 ( .A1(n1013), .A2(n1017), .ZN(n1187) );
  NAND2_X1 U1171 ( .A1(n895), .A2(n894), .ZN(n1252) );
  FA_X1 U1172 ( .A(\intadd_23/SUM[2] ), .B(\intadd_22/SUM[1] ), .CI(
        \intadd_35/n1 ), .CO(n896), .S(n895) );
  NAND2_X1 U1173 ( .A1(\intadd_23/SUM[3] ), .A2(n896), .ZN(n1249) );
  NAND2_X1 U1174 ( .A1(n1252), .A2(n1249), .ZN(n1028) );
  NOR2_X1 U1175 ( .A1(n1187), .A2(n1028), .ZN(n1030) );
  OAI21_X1 U1176 ( .B1(\intadd_23/SUM[2] ), .B2(\intadd_35/n1 ), .A(
        \intadd_22/SUM[1] ), .ZN(n898) );
  AOI21_X1 U1177 ( .B1(\intadd_35/n1 ), .B2(\intadd_23/SUM[2] ), .A(
        \intadd_23/SUM[3] ), .ZN(n897) );
  NAND2_X1 U1178 ( .A1(n898), .A2(n897), .ZN(n1248) );
  OAI21_X1 U1179 ( .B1(\intadd_23/n1 ), .B2(\intadd_22/SUM[3] ), .A(n1248), 
        .ZN(n1188) );
  NOR2_X1 U1180 ( .A1(n1030), .A2(n1188), .ZN(n1225) );
  NOR2_X1 U1181 ( .A1(n900), .A2(n899), .ZN(n1033) );
  NAND2_X1 U1182 ( .A1(\intadd_7/SUM[2] ), .A2(n925), .ZN(n901) );
  NAND2_X1 U1183 ( .A1(n901), .A2(n902), .ZN(n1244) );
  FA_X1 U1184 ( .A(\intadd_6/SUM[1] ), .B(\intadd_33/n1 ), .CI(n1001), .CO(
        n946), .S(n397) );
  AOI21_X1 U1185 ( .B1(\intadd_10/n1 ), .B2(n1244), .A(n1243), .ZN(n924) );
  NAND2_X1 U1186 ( .A1(\intadd_7/SUM[2] ), .A2(n903), .ZN(n923) );
  AOI22_X1 U1187 ( .A1(\intadd_10/n1 ), .A2(\intadd_11/B[3] ), .B1(
        \intadd_9/n1 ), .B2(\intadd_10/SUM[4] ), .ZN(n921) );
  NAND2_X1 U1188 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
  NOR2_X1 U1189 ( .A1(\intadd_31/n1 ), .A2(\intadd_9/SUM[3] ), .ZN(n907) );
  OAI221_X1 U1190 ( .B1(\intadd_31/n1 ), .B2(\intadd_10/SUM[2] ), .C1(
        \intadd_31/n1 ), .C2(\intadd_21/n1 ), .A(\intadd_11/A[1] ), .ZN(n906)
         );
  NOR4_X1 U1191 ( .A1(\intadd_31/n1 ), .A2(\intadd_10/SUM[2] ), .A3(
        \intadd_21/n1 ), .A4(\intadd_9/SUM[3] ), .ZN(n905) );
  OAI22_X1 U1192 ( .A1(n907), .A2(n906), .B1(n905), .B2(n904), .ZN(n919) );
  INV_X2 U1193 ( .A(\intadd_30/n1 ), .ZN(n916) );
  NOR2_X1 U1194 ( .A1(\intadd_31/SUM[2] ), .A2(n916), .ZN(n1209) );
  AOI21_X1 U1195 ( .B1(n910), .B2(n909), .A(n908), .ZN(n911) );
  AOI22_X1 U1196 ( .A1(n912), .A2(n911), .B1(\intadd_20/n1 ), .B2(
        \intadd_19/SUM[3] ), .ZN(n914) );
  OAI22_X1 U1197 ( .A1(\intadd_20/n1 ), .A2(\intadd_19/SUM[3] ), .B1(
        \intadd_19/n1 ), .B2(n1212), .ZN(n913) );
  NOR2_X1 U1198 ( .A1(n914), .A2(n913), .ZN(n915) );
  AOI21_X1 U1199 ( .B1(\intadd_19/n1 ), .B2(n1212), .A(n915), .ZN(n1058) );
  AOI22_X1 U1200 ( .A1(\intadd_9/SUM[4] ), .A2(\intadd_11/A[1] ), .B1(
        \intadd_11/B[0] ), .B2(\intadd_31/n1 ), .ZN(n917) );
  NAND2_X1 U1201 ( .A1(\intadd_31/SUM[2] ), .A2(n916), .ZN(n1208) );
  OAI211_X1 U1202 ( .C1(n1209), .C2(n1058), .A(n917), .B(n1208), .ZN(n918) );
  OAI211_X1 U1203 ( .C1(\intadd_9/n1 ), .C2(\intadd_10/SUM[4] ), .A(n919), .B(
        n918), .ZN(n920) );
  AND3_X1 U1204 ( .A1(n921), .A2(n1242), .A3(n920), .ZN(n922) );
  AOI21_X1 U1205 ( .B1(n924), .B2(n923), .A(n922), .ZN(n1075) );
  OR3_X1 U1206 ( .A1(\intadd_7/SUM[2] ), .A2(\intadd_10/n1 ), .A3(n925), .ZN(
        n1074) );
  FA_X1 U1207 ( .A(\intadd_25/SUM[1] ), .B(n926), .CI(\intadd_3/SUM[1] ), .CO(
        \intadd_4/B[3] ), .S(n953) );
  AOI222_X1 U1208 ( .A1(n953), .A2(\intadd_15/n1 ), .B1(n953), .B2(
        \intadd_17/SUM[3] ), .C1(\intadd_15/n1 ), .C2(\intadd_17/SUM[3] ), 
        .ZN(n971) );
  NOR2_X1 U1209 ( .A1(\intadd_4/SUM[3] ), .A2(\intadd_25/SUM[2] ), .ZN(n952)
         );
  AOI21_X1 U1210 ( .B1(\intadd_25/SUM[2] ), .B2(\intadd_4/SUM[3] ), .A(n952), 
        .ZN(n927) );
  XNOR2_X1 U1211 ( .A(\intadd_17/n1 ), .B(n927), .ZN(n970) );
  NOR2_X1 U1212 ( .A1(n971), .A2(n970), .ZN(n1082) );
  FA_X1 U1213 ( .A(n930), .B(n929), .CI(n928), .CO(\intadd_5/B[3] ), .S(n957)
         );
  FA_X1 U1214 ( .A(n933), .B(n932), .CI(n931), .CO(n937), .S(\intadd_6/A[4] )
         );
  AOI22_X1 U1215 ( .A1(\intadd_6/n1 ), .A2(n954), .B1(\intadd_7/n1 ), .B2(
        \intadd_6/SUM[4] ), .ZN(n1008) );
  AOI21_X1 U1216 ( .B1(\intadd_16/n1 ), .B2(n956), .A(n957), .ZN(n934) );
  FA_X1 U1217 ( .A(n936), .B(n935), .CI(\intadd_17/SUM[1] ), .CO(
        \intadd_15/B[3] ), .S(n941) );
  FA_X1 U1218 ( .A(\intadd_27/n1 ), .B(\intadd_5/SUM[2] ), .CI(n937), .CO(n942), .S(n956) );
  AOI221_X1 U1219 ( .B1(\intadd_27/n1 ), .B2(n938), .C1(\intadd_5/SUM[2] ), 
        .C2(n937), .A(n941), .ZN(n945) );
  AOI21_X1 U1220 ( .B1(n941), .B2(n942), .A(n945), .ZN(n939) );
  XOR2_X1 U1221 ( .A(\intadd_5/SUM[3] ), .B(n939), .Z(n959) );
  OAI211_X1 U1222 ( .C1(n956), .C2(\intadd_16/n1 ), .A(n940), .B(n959), .ZN(
        n995) );
  NAND2_X1 U1223 ( .A1(n942), .A2(n941), .ZN(n943) );
  OAI21_X1 U1224 ( .B1(n945), .B2(n944), .A(n943), .ZN(n961) );
  NAND2_X1 U1225 ( .A1(\intadd_5/SUM[4] ), .A2(n961), .ZN(n1196) );
  NAND2_X1 U1226 ( .A1(\intadd_3/SUM[4] ), .A2(\intadd_4/n1 ), .ZN(n1181) );
  AOI21_X1 U1227 ( .B1(\intadd_25/SUM[2] ), .B2(\intadd_4/SUM[3] ), .A(
        \intadd_17/n1 ), .ZN(n951) );
  NOR2_X1 U1228 ( .A1(n952), .A2(n974), .ZN(n1255) );
  NAND2_X1 U1229 ( .A1(n996), .A2(\intadd_5/n1 ), .ZN(n997) );
  NOR3_X1 U1230 ( .A1(n972), .A2(n1255), .A3(n1084), .ZN(n963) );
  AND3_X1 U1231 ( .A1(n995), .A2(n1196), .A3(n963), .ZN(n947) );
  FA_X1 U1232 ( .A(\intadd_7/SUM[3] ), .B(n946), .CI(\intadd_6/SUM[2] ), .CO(
        n1003), .S(n1243) );
  NAND2_X1 U1233 ( .A1(n1003), .A2(\intadd_7/SUM[4] ), .ZN(n1002) );
  NAND3_X1 U1234 ( .A1(n1008), .A2(n947), .A3(n1002), .ZN(n948) );
  AOI211_X1 U1235 ( .C1(n1075), .C2(n1074), .A(n1082), .B(n948), .ZN(n1022) );
  AOI21_X1 U1236 ( .B1(\intadd_13/B[3] ), .B2(\intadd_13/A[3] ), .A(
        \intadd_14/SUM[3] ), .ZN(n949) );
  NAND2_X1 U1237 ( .A1(\intadd_13/SUM[3] ), .A2(\intadd_2/n1 ), .ZN(n1066) );
  NAND2_X1 U1238 ( .A1(\intadd_14/SUM[3] ), .A2(\intadd_13/n1 ), .ZN(n1062) );
  OAI21_X1 U1239 ( .B1(n949), .B2(n1066), .A(n1062), .ZN(n1130) );
  NAND2_X1 U1240 ( .A1(\intadd_3/n1 ), .A2(\intadd_1/SUM[4] ), .ZN(n1180) );
  NAND2_X1 U1241 ( .A1(\intadd_2/SUM[4] ), .A2(\intadd_1/n1 ), .ZN(n1019) );
  NAND2_X1 U1242 ( .A1(n1180), .A2(n1019), .ZN(n1059) );
  NOR2_X1 U1243 ( .A1(n1130), .A2(n1059), .ZN(n979) );
  OAI21_X1 U1244 ( .B1(n952), .B2(n951), .A(n950), .ZN(n1010) );
  OAI21_X1 U1245 ( .B1(\intadd_3/SUM[4] ), .B2(\intadd_4/n1 ), .A(n1010), .ZN(
        n1183) );
  FA_X1 U1246 ( .A(n953), .B(\intadd_15/n1 ), .CI(\intadd_17/SUM[3] ), .CO(
        n967), .S(n996) );
  NAND2_X1 U1247 ( .A1(n995), .A2(n1196), .ZN(n1083) );
  NOR2_X1 U1248 ( .A1(n1003), .A2(\intadd_7/SUM[4] ), .ZN(n1072) );
  NOR2_X1 U1249 ( .A1(\intadd_7/n1 ), .A2(\intadd_6/SUM[4] ), .ZN(n955) );
  NAND2_X1 U1250 ( .A1(\intadd_6/n1 ), .A2(n954), .ZN(n1089) );
  NOR2_X1 U1251 ( .A1(\intadd_6/n1 ), .A2(n954), .ZN(n1090) );
  AOI21_X1 U1252 ( .B1(n955), .B2(n1089), .A(n1090), .ZN(n1009) );
  FA_X1 U1253 ( .A(n957), .B(\intadd_16/n1 ), .CI(n956), .CO(n958), .S(n954)
         );
  NOR2_X1 U1254 ( .A1(n959), .A2(n958), .ZN(n1177) );
  NAND2_X1 U1255 ( .A1(n1009), .A2(n960), .ZN(n1258) );
  AOI21_X1 U1256 ( .B1(n1072), .B2(n1008), .A(n1258), .ZN(n962) );
  NOR2_X1 U1257 ( .A1(\intadd_5/SUM[4] ), .A2(n961), .ZN(n1198) );
  NOR2_X1 U1258 ( .A1(n996), .A2(\intadd_5/n1 ), .ZN(n1078) );
  NOR2_X1 U1259 ( .A1(n1198), .A2(n1078), .ZN(n1257) );
  OAI21_X1 U1260 ( .B1(n1083), .B2(n962), .A(n1257), .ZN(n964) );
  NAND2_X1 U1261 ( .A1(n964), .A2(n963), .ZN(n965) );
  AOI21_X1 U1262 ( .B1(n967), .B2(n966), .A(n965), .ZN(n969) );
  NOR2_X1 U1263 ( .A1(\intadd_3/n1 ), .A2(\intadd_1/SUM[4] ), .ZN(n968) );
  AOI211_X1 U1264 ( .C1(n1181), .C2(n1183), .A(n969), .B(n968), .ZN(n1020) );
  NAND2_X1 U1265 ( .A1(n971), .A2(n970), .ZN(n1265) );
  NOR2_X1 U1266 ( .A1(n972), .A2(n1265), .ZN(n1024) );
  NOR2_X1 U1267 ( .A1(\intadd_14/SUM[3] ), .A2(\intadd_13/n1 ), .ZN(n1061) );
  NOR2_X1 U1268 ( .A1(\intadd_2/SUM[4] ), .A2(\intadd_1/n1 ), .ZN(n1202) );
  OAI21_X1 U1269 ( .B1(\intadd_13/SUM[3] ), .B2(\intadd_2/n1 ), .A(n1065), 
        .ZN(n1067) );
  NOR2_X1 U1270 ( .A1(n1061), .A2(n1067), .ZN(n1133) );
  AOI21_X1 U1271 ( .B1(n1024), .B2(n974), .A(n973), .ZN(n977) );
  AOI21_X1 U1272 ( .B1(n1133), .B2(n1059), .A(n1130), .ZN(n975) );
  AOI21_X1 U1273 ( .B1(n1020), .B2(n977), .A(n976), .ZN(n978) );
  AOI21_X1 U1274 ( .B1(n1022), .B2(n979), .A(n978), .ZN(n1226) );
  NOR3_X1 U1275 ( .A1(n1033), .A2(n1226), .A3(n1028), .ZN(n980) );
  NAND2_X1 U1276 ( .A1(\intadd_23/n1 ), .A2(\intadd_22/SUM[3] ), .ZN(n1119) );
  OAI21_X1 U1277 ( .B1(n981), .B2(n980), .A(n1119), .ZN(n994) );
  FA_X1 U1278 ( .A(n984), .B(n983), .CI(n982), .CO(n1112), .S(n990) );
  NOR2_X1 U1279 ( .A1(n575), .A2(n824), .ZN(n987) );
  OAI21_X1 U1280 ( .B1(n987), .B2(n986), .A(n985), .ZN(n1111) );
  AOI22_X1 U1281 ( .A1(b[19]), .A2(n1150), .B1(n1108), .B2(n1106), .ZN(n988)
         );
  AOI221_X1 U1282 ( .B1(n1139), .B2(b[20]), .C1(n1147), .C2(n1098), .A(n988), 
        .ZN(n1110) );
  FA_X1 U1283 ( .A(n991), .B(n990), .CI(n989), .CO(n1121), .S(\intadd_22/B[3] ) );
  NAND2_X1 U1284 ( .A1(\intadd_22/n1 ), .A2(n992), .ZN(n1120) );
  NOR2_X1 U1285 ( .A1(\intadd_22/n1 ), .A2(n992), .ZN(n1228) );
  INV_X1 U1286 ( .A(n1228), .ZN(n1190) );
  NAND2_X1 U1287 ( .A1(n1120), .A2(n1190), .ZN(n993) );
  XNOR2_X1 U1288 ( .A(n994), .B(n993), .ZN(\d[42]_BAR ) );
  AOI21_X1 U1289 ( .B1(\intadd_5/B[4] ), .B2(\intadd_5/A[4] ), .A(n996), .ZN(
        n998) );
  OAI21_X1 U1290 ( .B1(n998), .B2(n1196), .A(n997), .ZN(n999) );
  AOI21_X1 U1291 ( .B1(n1257), .B2(n1194), .A(n999), .ZN(n1261) );
  NOR4_X1 U1292 ( .A1(\intadd_10/n1 ), .A2(\intadd_7/SUM[2] ), .A3(
        \intadd_7/SUM[4] ), .A4(n1000), .ZN(n1006) );
  NAND3_X1 U1293 ( .A1(\intadd_6/SUM[1] ), .A2(\intadd_33/n1 ), .A3(n1001), 
        .ZN(n1005) );
  OAI22_X1 U1294 ( .A1(n1003), .A2(n1074), .B1(n1075), .B2(n1073), .ZN(n1004)
         );
  AOI211_X1 U1295 ( .C1(n1006), .C2(n1005), .A(n1072), .B(n1004), .ZN(n1092)
         );
  NAND2_X1 U1296 ( .A1(n1008), .A2(n1007), .ZN(n1262) );
  NAND2_X1 U1297 ( .A1(n1009), .A2(n1262), .ZN(n1176) );
  NOR2_X1 U1298 ( .A1(n1177), .A2(n1176), .ZN(n1195) );
  NAND2_X1 U1299 ( .A1(n1257), .A2(n1195), .ZN(n1264) );
  NAND2_X1 U1300 ( .A1(n1261), .A2(n1264), .ZN(n1088) );
  AOI211_X1 U1301 ( .C1(n1265), .C2(n1088), .A(n1082), .B(n1255), .ZN(n1182)
         );
  NOR2_X1 U1302 ( .A1(n1182), .A2(n1256), .ZN(n1012) );
  OAI21_X1 U1303 ( .B1(\intadd_3/SUM[4] ), .B2(\intadd_4/n1 ), .A(n1181), .ZN(
        n1011) );
  XNOR2_X1 U1304 ( .A(n1012), .B(n1011), .ZN(\d[33]_BAR ) );
  INV_X1 U1305 ( .A(n1013), .ZN(n1032) );
  NAND2_X1 U1306 ( .A1(n1252), .A2(n1032), .ZN(n1016) );
  OAI21_X1 U1307 ( .B1(n1017), .B2(n1014), .A(n1029), .ZN(n1015) );
  XNOR2_X1 U1308 ( .A(n1016), .B(n1015), .ZN(\d[39]_BAR ) );
  NOR2_X1 U1309 ( .A1(n1033), .A2(n1017), .ZN(n1018) );
  XOR2_X1 U1310 ( .A(n1018), .B(n1226), .Z(\d[38]_BAR ) );
  NAND2_X1 U1311 ( .A1(n1065), .A2(n1019), .ZN(n1027) );
  INV_X1 U1312 ( .A(n1180), .ZN(n1025) );
  AOI211_X1 U1313 ( .C1(n1024), .C2(n1023), .A(n1022), .B(n1021), .ZN(n1060)
         );
  NOR2_X1 U1314 ( .A1(n1025), .A2(n1060), .ZN(n1026) );
  XNOR2_X1 U1315 ( .A(n1027), .B(n1026), .ZN(\d[35] ) );
  OAI21_X1 U1316 ( .B1(\intadd_23/n1 ), .B2(\intadd_22/SUM[3] ), .A(n1119), 
        .ZN(n1039) );
  NAND2_X1 U1317 ( .A1(n1034), .A2(n1029), .ZN(n1129) );
  INV_X1 U1318 ( .A(n1030), .ZN(n1031) );
  OAI211_X1 U1319 ( .C1(n1226), .C2(n1129), .A(n1248), .B(n1031), .ZN(n1038)
         );
  NAND2_X1 U1320 ( .A1(n1033), .A2(n1032), .ZN(n1250) );
  NAND2_X1 U1321 ( .A1(n1034), .A2(n1250), .ZN(n1224) );
  AOI21_X1 U1322 ( .B1(n1226), .B2(n1187), .A(n1224), .ZN(n1036) );
  NOR3_X1 U1323 ( .A1(n1039), .A2(n1036), .A3(n1035), .ZN(n1037) );
  AOI21_X1 U1324 ( .B1(n1039), .B2(n1038), .A(n1037), .ZN(\d[41]_BAR ) );
  XOR2_X1 U1325 ( .A(n1041), .B(n1040), .Z(\d[2] ) );
  INV_X1 U1326 ( .A(n1042), .ZN(n1044) );
  NOR2_X1 U1327 ( .A1(n1044), .A2(n1043), .ZN(n1049) );
  AOI22_X1 U1328 ( .A1(n1047), .A2(\intadd_26/SUM[0] ), .B1(n1046), .B2(n1045), 
        .ZN(n1048) );
  XNOR2_X1 U1329 ( .A(n1049), .B(n1048), .ZN(\d[5]_BAR ) );
  OAI222_X1 U1330 ( .A1(\intadd_26/n1 ), .A2(n1051), .B1(\intadd_26/n1 ), .B2(
        n1054), .C1(n1050), .C2(n1055), .ZN(\d[8]_BAR ) );
  AOI21_X1 U1331 ( .B1(n1053), .B2(\intadd_8/SUM[1] ), .A(n1052), .ZN(n1057)
         );
  NAND2_X1 U1332 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  XNOR2_X1 U1333 ( .A(n1057), .B(n1056), .ZN(\d[9]_BAR ) );
  AOI21_X1 U1334 ( .B1(n1058), .B2(n1208), .A(n1209), .ZN(\intadd_11/CI ) );
  NOR2_X1 U1335 ( .A1(n1060), .A2(n1059), .ZN(n1201) );
  NAND2_X1 U1336 ( .A1(n1201), .A2(n1066), .ZN(n1064) );
  NAND2_X1 U1337 ( .A1(n1063), .A2(n1062), .ZN(n1069) );
  NAND2_X1 U1338 ( .A1(n1064), .A2(n1069), .ZN(n1071) );
  INV_X1 U1339 ( .A(n1066), .ZN(n1203) );
  OAI22_X1 U1340 ( .A1(\intadd_13/SUM[3] ), .A2(\intadd_2/n1 ), .B1(n1203), 
        .B2(n1065), .ZN(n1070) );
  OAI21_X1 U1341 ( .B1(n1201), .B2(n1067), .A(n1066), .ZN(n1068) );
  OAI22_X1 U1342 ( .A1(n1071), .A2(n1070), .B1(n1069), .B2(n1068), .ZN(
        \d[37]_BAR ) );
  NOR2_X1 U1343 ( .A1(n1073), .A2(n1072), .ZN(n1077) );
  NAND2_X1 U1344 ( .A1(n1075), .A2(n1074), .ZN(n1076) );
  XOR2_X1 U1345 ( .A(n1077), .B(n1076), .Z(\d[25] ) );
  NOR2_X1 U1346 ( .A1(n1078), .A2(n1084), .ZN(n1081) );
  NOR2_X1 U1347 ( .A1(n1195), .A2(n1083), .ZN(n1079) );
  NOR2_X1 U1348 ( .A1(n1198), .A2(n1079), .ZN(n1080) );
  XNOR2_X1 U1349 ( .A(n1081), .B(n1080), .ZN(\d[30] ) );
  INV_X1 U1350 ( .A(n1082), .ZN(n1260) );
  NAND2_X1 U1351 ( .A1(n1260), .A2(n1265), .ZN(n1087) );
  OAI21_X1 U1352 ( .B1(n1195), .B2(n1083), .A(n1257), .ZN(n1086) );
  NOR2_X1 U1353 ( .A1(n1087), .A2(n1084), .ZN(n1085) );
  AOI22_X1 U1354 ( .A1(n1088), .A2(n1087), .B1(n1086), .B2(n1085), .ZN(\d[31] ) );
  NOR2_X1 U1355 ( .A1(n1091), .A2(n1090), .ZN(n1094) );
  FA_X1 U1356 ( .A(\intadd_6/SUM[4] ), .B(\intadd_7/n1 ), .CI(n1092), .CO(
        n1093), .S(\d[26]_BAR ) );
  XOR2_X1 U1357 ( .A(n1094), .B(n1093), .Z(\d[27]_BAR ) );
  NOR2_X1 U1358 ( .A1(a[19]), .A2(n1095), .ZN(n1097) );
  AOI221_X1 U1359 ( .B1(n1101), .B2(b[23]), .C1(n1097), .C2(n1163), .A(n1096), 
        .ZN(n1146) );
  NOR2_X1 U1360 ( .A1(n1105), .A2(n1098), .ZN(n1153) );
  AOI22_X1 U1361 ( .A1(b[21]), .A2(n1150), .B1(n1108), .B2(n878), .ZN(n1099)
         );
  AOI221_X1 U1362 ( .B1(n1139), .B2(b[22]), .C1(n1147), .C2(n1140), .A(n1099), 
        .ZN(n1145) );
  NOR2_X1 U1363 ( .A1(n1114), .A2(n1106), .ZN(n1107) );
  AOI22_X1 U1364 ( .A1(b[22]), .A2(n1101), .B1(n1100), .B2(n1140), .ZN(n1102)
         );
  OAI221_X1 U1365 ( .B1(b[23]), .B2(n1104), .C1(n1151), .C2(n1103), .A(n1102), 
        .ZN(n1115) );
  AOI21_X1 U1366 ( .B1(n1114), .B2(n1106), .A(n1105), .ZN(n1113) );
  OAI21_X1 U1367 ( .B1(n1107), .B2(n1115), .A(n1113), .ZN(\intadd_12/B[2] ) );
  AOI22_X1 U1368 ( .A1(b[20]), .A2(n1150), .B1(n1108), .B2(n1098), .ZN(n1109)
         );
  AOI221_X1 U1369 ( .B1(n1139), .B2(b[21]), .C1(n1147), .C2(n878), .A(n1109), 
        .ZN(\intadd_12/B[1] ) );
  FA_X1 U1370 ( .A(n1112), .B(n1111), .CI(n1110), .CO(n1126), .S(n1122) );
  OAI21_X1 U1371 ( .B1(n1106), .B2(n1114), .A(n1113), .ZN(n1116) );
  XOR2_X1 U1372 ( .A(n1116), .B(n1115), .Z(n1125) );
  NAND2_X1 U1373 ( .A1(\intadd_12/SUM[2] ), .A2(n1117), .ZN(n1222) );
  AND2_X1 U1374 ( .A1(\intadd_12/SUM[0] ), .A2(n1122), .ZN(n1118) );
  FA_X1 U1375 ( .A(n1126), .B(\intadd_12/SUM[1] ), .CI(n1125), .CO(n1117), .S(
        n1124) );
  OAI221_X1 U1376 ( .B1(\intadd_12/SUM[0] ), .B2(n1122), .C1(n1121), .C2(n1118), .A(n1124), .ZN(n1229) );
  NAND2_X1 U1377 ( .A1(n1222), .A2(n1229), .ZN(n1231) );
  NAND2_X1 U1378 ( .A1(n1120), .A2(n1119), .ZN(n1223) );
  FA_X1 U1379 ( .A(n1122), .B(\intadd_12/SUM[0] ), .CI(n1121), .CO(n1123), .S(
        n992) );
  NOR2_X1 U1380 ( .A1(n1124), .A2(n1123), .ZN(n1227) );
  NOR2_X1 U1381 ( .A1(n1227), .A2(n1228), .ZN(n1233) );
  OAI21_X1 U1382 ( .B1(n1225), .B2(n1223), .A(n1233), .ZN(n1136) );
  OAI21_X1 U1383 ( .B1(\intadd_12/SUM[1] ), .B2(n1126), .A(n1125), .ZN(n1128)
         );
  AOI21_X1 U1384 ( .B1(n1126), .B2(\intadd_12/SUM[1] ), .A(\intadd_12/SUM[2] ), 
        .ZN(n1127) );
  NAND2_X1 U1385 ( .A1(n1128), .A2(n1127), .ZN(n1234) );
  INV_X1 U1386 ( .A(n1234), .ZN(n1135) );
  OR4_X1 U1387 ( .A1(n1130), .A2(n1223), .A3(n1231), .A4(n1129), .ZN(n1131) );
  AOI21_X1 U1388 ( .B1(n1133), .B2(n1132), .A(n1131), .ZN(n1134) );
  AOI211_X1 U1389 ( .C1(n1137), .C2(n1136), .A(n1135), .B(n1134), .ZN(
        \intadd_12/B[3] ) );
  AOI22_X1 U1390 ( .A1(b[23]), .A2(n1139), .B1(b[22]), .B2(n1138), .ZN(n1142)
         );
  AOI22_X1 U1391 ( .A1(n1141), .A2(n1140), .B1(n1147), .B2(n1151), .ZN(n1157)
         );
  NAND2_X1 U1392 ( .A1(n1142), .A2(n1157), .ZN(n1144) );
  NOR2_X1 U1393 ( .A1(n1153), .A2(b[21]), .ZN(n1154) );
  AOI211_X1 U1394 ( .C1(b[21]), .C2(b[20]), .A(n1154), .B(n1105), .ZN(n1143)
         );
  XNOR2_X1 U1395 ( .A(n1144), .B(n1143), .ZN(n1160) );
  FA_X1 U1396 ( .A(n1146), .B(n1153), .CI(n1145), .CO(n1159), .S(
        \intadd_12/A[2] ) );
  NOR2_X1 U1397 ( .A1(a[22]), .A2(n1105), .ZN(n1148) );
  AOI21_X1 U1398 ( .B1(n1148), .B2(n1151), .A(n1147), .ZN(n1155) );
  OAI211_X1 U1399 ( .C1(n1153), .C2(b[21]), .A(n1148), .B(n1140), .ZN(n1149)
         );
  OAI211_X1 U1400 ( .C1(n1151), .C2(n1150), .A(n1155), .B(n1149), .ZN(n1152)
         );
  AOI21_X1 U1401 ( .B1(n1153), .B2(b[21]), .A(n1152), .ZN(n1166) );
  NAND2_X1 U1402 ( .A1(n1153), .A2(b[21]), .ZN(n1156) );
  AOI211_X1 U1403 ( .C1(n1157), .C2(n1156), .A(n1155), .B(n1154), .ZN(n1167)
         );
  NOR2_X1 U1404 ( .A1(n1166), .A2(n1167), .ZN(n1158) );
  NAND2_X1 U1405 ( .A1(b[22]), .A2(a[23]), .ZN(n1165) );
  XNOR2_X1 U1406 ( .A(n1158), .B(n1165), .ZN(n1220) );
  FA_X1 U1407 ( .A(n1161), .B(n1160), .CI(n1159), .CO(n1221), .S(
        \intadd_12/A[3] ) );
  AOI21_X1 U1408 ( .B1(n1220), .B2(n1221), .A(\intadd_12/n1 ), .ZN(n1175) );
  OR2_X1 U1409 ( .A1(n1220), .A2(n1221), .ZN(n1171) );
  AOI221_X1 U1410 ( .B1(b[23]), .B2(n1164), .C1(n1163), .C2(n1162), .A(n1105), 
        .ZN(n1170) );
  INV_X1 U1411 ( .A(n1165), .ZN(n1168) );
  AOI22_X1 U1412 ( .A1(n1168), .A2(n1167), .B1(n1166), .B2(n1165), .ZN(n1169)
         );
  XNOR2_X1 U1413 ( .A(n1170), .B(n1169), .ZN(n1172) );
  NAND2_X1 U1414 ( .A1(n1171), .A2(n1172), .ZN(n1174) );
  OAI22_X1 U1415 ( .A1(n1175), .A2(n1174), .B1(n1173), .B2(n1172), .ZN(\d[47] ) );
  OAI21_X1 U1416 ( .B1(n1194), .B2(n1177), .A(n1176), .ZN(n1178) );
  OAI21_X1 U1417 ( .B1(n1194), .B2(n1179), .A(n1178), .ZN(\d[28] ) );
  OAI21_X1 U1418 ( .B1(\intadd_3/n1 ), .B2(\intadd_1/SUM[4] ), .A(n1180), .ZN(
        n1185) );
  OAI21_X1 U1419 ( .B1(n1183), .B2(n1182), .A(n1181), .ZN(n1184) );
  XOR2_X1 U1420 ( .A(n1185), .B(n1184), .Z(\d[34] ) );
  INV_X1 U1421 ( .A(n1227), .ZN(n1186) );
  NAND2_X1 U1422 ( .A1(n1229), .A2(n1186), .ZN(n1193) );
  INV_X1 U1423 ( .A(n1224), .ZN(n1189) );
  NAND2_X1 U1424 ( .A1(n1187), .A2(n1226), .ZN(n1251) );
  AOI21_X1 U1425 ( .B1(n1189), .B2(n1251), .A(n1188), .ZN(n1191) );
  OAI21_X1 U1426 ( .B1(n1191), .B2(n1223), .A(n1190), .ZN(n1192) );
  XNOR2_X1 U1427 ( .A(n1193), .B(n1192), .ZN(\d[43] ) );
  NOR2_X1 U1428 ( .A1(n1195), .A2(n1194), .ZN(n1200) );
  INV_X1 U1429 ( .A(n1196), .ZN(n1197) );
  NOR2_X1 U1430 ( .A1(n1198), .A2(n1197), .ZN(n1199) );
  XOR2_X1 U1431 ( .A(n1200), .B(n1199), .Z(\d[29] ) );
  NOR2_X1 U1432 ( .A1(n1202), .A2(n1201), .ZN(n1206) );
  NOR2_X1 U1433 ( .A1(\intadd_13/SUM[3] ), .A2(\intadd_2/n1 ), .ZN(n1204) );
  NOR2_X1 U1434 ( .A1(n1204), .A2(n1203), .ZN(n1205) );
  XOR2_X1 U1435 ( .A(n1206), .B(n1205), .Z(\d[36]_BAR ) );
  FA_X1 U1436 ( .A(\intadd_20/n1 ), .B(\intadd_19/SUM[3] ), .CI(n1207), .CO(
        n1211), .S(\d[17]_BAR ) );
  INV_X1 U1437 ( .A(n1208), .ZN(n1210) );
  NOR2_X1 U1438 ( .A1(n1210), .A2(n1209), .ZN(n1214) );
  FA_X1 U1439 ( .A(\intadd_19/n1 ), .B(n1212), .CI(n1211), .CO(n1213), .S(n13)
         );
  XNOR2_X1 U1440 ( .A(n1214), .B(n1213), .ZN(\d[19] ) );
  AOI21_X1 U1441 ( .B1(\intadd_20/SUM[3] ), .B2(n1216), .A(n1215), .ZN(n1218)
         );
  XNOR2_X1 U1442 ( .A(n1218), .B(n1217), .ZN(\d[16] ) );
  FA_X1 U1443 ( .A(\intadd_18/n1 ), .B(\intadd_0/n1 ), .CI(n1219), .CO(n1217), 
        .S(\d[15]_BAR ) );
  FA_X1 U1444 ( .A(\intadd_12/n1 ), .B(n1221), .CI(n1220), .CO(n1173), .S(
        \d[46]_BAR ) );
  NAND2_X1 U1445 ( .A1(n1234), .A2(n1222), .ZN(n1237) );
  AOI221_X1 U1446 ( .B1(n1226), .B2(n1225), .C1(n1224), .C2(n1225), .A(n1223), 
        .ZN(n1230) );
  AOI221_X1 U1447 ( .B1(n1230), .B2(n1229), .C1(n1228), .C2(n1229), .A(n1227), 
        .ZN(n1236) );
  AOI21_X1 U1448 ( .B1(n1233), .B2(n1232), .A(n1231), .ZN(n1235) );
  AOI22_X1 U1449 ( .A1(n1237), .A2(n1236), .B1(n1235), .B2(n1234), .ZN(\d[44] ) );
  NOR2_X1 U1450 ( .A1(n1239), .A2(n1238), .ZN(n1241) );
  NAND2_X1 U1451 ( .A1(b[1]), .A2(a[0]), .ZN(n1240) );
  XNOR2_X1 U1452 ( .A(n1241), .B(n1240), .ZN(\d[1] ) );
  OAI21_X1 U1453 ( .B1(n1244), .B2(n1243), .A(n1242), .ZN(n1245) );
  XNOR2_X1 U1454 ( .A(n1245), .B(\intadd_11/n1 ), .ZN(\d[24]_BAR ) );
  NOR2_X1 U1455 ( .A1(n1247), .A2(n1246), .ZN(\d[0] ) );
  NAND2_X1 U1456 ( .A1(n1249), .A2(n1248), .ZN(n1254) );
  NAND3_X1 U1457 ( .A1(n1252), .A2(n1251), .A3(n1250), .ZN(n1253) );
  XOR2_X1 U1458 ( .A(n1254), .B(n1253), .Z(\d[40] ) );
  NOR2_X1 U1459 ( .A1(n1256), .A2(n1255), .ZN(n1269) );
  NAND2_X1 U1460 ( .A1(n1269), .A2(n1265), .ZN(n1272) );
  INV_X1 U1461 ( .A(n1257), .ZN(n1259) );
  NOR2_X1 U1462 ( .A1(n1259), .A2(n1258), .ZN(n1263) );
  NAND2_X1 U1463 ( .A1(n1261), .A2(n1260), .ZN(n1267) );
  AOI21_X1 U1464 ( .B1(n1263), .B2(n1262), .A(n1267), .ZN(n1271) );
  OAI21_X1 U1465 ( .B1(n1267), .B2(n1266), .A(n1265), .ZN(n1268) );
  OAI22_X1 U1466 ( .A1(n1272), .A2(n1271), .B1(n1270), .B2(n1269), .ZN(\d[32] ) );
  FA_X1 U1467 ( .A(n1275), .B(n1274), .CI(n1273), .CO(n1281), .S(\d[3]_BAR )
         );
  AOI22_X1 U1468 ( .A1(n1279), .A2(n1278), .B1(n1277), .B2(n1276), .ZN(n1280)
         );
  XNOR2_X1 U1469 ( .A(n1281), .B(n1280), .ZN(\d[4]_BAR ) );
  AND2_X1 U6 ( .A1(n497), .A2(a[11]), .ZN(n793) );
  INV_X1 U7 ( .A(a[23]), .ZN(n1105) );
endmodule



    module conf_int_mul__noFF__arch_agnos__w_wrapper_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 ( 
        clk, rst, a, b, d__acc, acc__sel, \d[63] , \d[62] , \d[61] , \d[60] , 
        \d[59] , \d[58] , \d[57] , \d[56] , \d[55] , \d[54] , \d[53] , \d[52] , 
        \d[51] , \d[50] , \d[49] , \d[48] , \d[47] , \d[46] , \d[45] , \d[44] , 
        \d[43] , \d[42] , \d[41] , \d[40] , \d[39] , \d[38] , \d[37] , \d[36] , 
        \d[35] , \d[34] , \d[33] , \d[32] , \d[31] , \d[30] , \d[29] , 
        \d[28]_BAR , \d[23] , \d[22] , \d[21] , \d[20] , \d[19] , \d[18] , 
        \d[17] , \d[16] , \d[15] , \d[14] , \d[13] , \d[12] , \d[11] , \d[10] , 
        \d[9] , \d[8] , \d[7] , \d[6] , \d[5] , \d[4] , \d[3] , \d[2] , \d[1] , 
        \d[0] , \d[27]_BAR , \d[26]_BAR , \d[25]_BAR , \d[24]_BAR  );
  input [23:0] a;
  input [23:0] b;
  input [63:0] d__acc;
  input clk, rst, acc__sel;
  output \d[63] , \d[62] , \d[61] , \d[60] , \d[59] , \d[58] , \d[57] ,
         \d[56] , \d[55] , \d[54] , \d[53] , \d[52] , \d[51] , \d[50] ,
         \d[49] , \d[48] , \d[47] , \d[46] , \d[45] , \d[44] , \d[43] ,
         \d[42] , \d[41] , \d[40] , \d[39] , \d[38] , \d[37] , \d[36] ,
         \d[35] , \d[34] , \d[33] , \d[32] , \d[31] , \d[30] , \d[29] ,
         \d[28]_BAR , \d[23] , \d[22] , \d[21] , \d[20] , \d[19] , \d[18] ,
         \d[17] , \d[16] , \d[15] , \d[14] , \d[13] , \d[12] , \d[11] ,
         \d[10] , \d[9] , \d[8] , \d[7] , \d[6] , \d[5] , \d[4] , \d[3] ,
         \d[2] , \d[1] , \d[0] , \d[27]_BAR , \d[26]_BAR , \d[25]_BAR ,
         \d[24]_BAR ;
  wire   n1, n2, n3, n4, n5, n6, n8, n10, n12, n14, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37;
  wire   [63:0] d;
  wire   [47:0] d__apx;
  assign \d[63]  = d[63];
  assign \d[62]  = d[62];
  assign \d[61]  = d[61];
  assign \d[60]  = d[60];
  assign \d[59]  = d[59];
  assign \d[58]  = d[58];
  assign \d[57]  = d[57];
  assign \d[56]  = d[56];
  assign \d[55]  = d[55];
  assign \d[54]  = d[54];
  assign \d[53]  = d[53];
  assign \d[52]  = d[52];
  assign \d[51]  = d[51];
  assign \d[50]  = d[50];
  assign \d[49]  = d[49];
  assign \d[48]  = d[48];
  assign \d[47]  = d[47];
  assign \d[46]  = d[46];
  assign \d[45]  = d[45];
  assign \d[44]  = d[44];
  assign \d[43]  = d[43];
  assign \d[42]  = d[42];
  assign \d[41]  = d[41];
  assign \d[40]  = d[40];
  assign \d[39]  = d[39];
  assign \d[38]  = d[38];
  assign \d[37]  = d[37];
  assign \d[36]  = d[36];
  assign \d[35]  = d[35];
  assign \d[34]  = d[34];
  assign \d[33]  = d[33];
  assign \d[32]  = d[32];
  assign \d[31]  = d[31];
  assign \d[30]  = d[30];
  assign \d[29]  = d[29];
  assign \d[23]  = d[23];
  assign \d[22]  = d[22];
  assign \d[21]  = d[21];
  assign \d[20]  = d[20];
  assign \d[18]  = d[18];
  assign \d[17]  = d[17];
  assign \d[16]  = d[16];
  assign \d[15]  = d[15];
  assign \d[14]  = d[14];
  assign \d[13]  = d[13];
  assign \d[12]  = d[12];
  assign \d[11]  = d[11];
  assign \d[10]  = d[10];
  assign \d[9]  = d[9];
  assign \d[8]  = d[8];
  assign \d[7]  = d[7];
  assign \d[6]  = d[6];
  assign \d[5]  = d[5];
  assign \d[4]  = d[4];
  assign \d[3]  = d[3];
  assign \d[2]  = d[2];
  assign \d[1]  = d[1];
  assign \d[0]  = d[0];

  INV_X1 U1 ( .A(d__apx[3]), .ZN(n2) );
  INV_X1 U2 ( .A(d__apx[6]), .ZN(n3) );
  INV_X1 U3 ( .A(d__apx[7]), .ZN(n4) );
  INV_X1 U4 ( .A(d__apx[12]), .ZN(n5) );
  LOGIC0_X1 U5 ( .Z(n1) );
  NOR2_X1 U6 ( .A1(d__apx[8]), .A2(acc__sel), .ZN(n6) );
  AOI21_X1 U7 ( .B1(d__acc[24]), .B2(acc__sel), .A(n6), .ZN(\d[24]_BAR ) );
  NOR2_X1 U8 ( .A1(d__apx[9]), .A2(acc__sel), .ZN(n8) );
  AOI21_X1 U9 ( .B1(d__acc[25]), .B2(acc__sel), .A(n8), .ZN(\d[25]_BAR ) );
  NOR2_X1 U10 ( .A1(d__apx[10]), .A2(acc__sel), .ZN(n10) );
  AOI21_X1 U11 ( .B1(d__acc[26]), .B2(acc__sel), .A(n10), .ZN(\d[26]_BAR ) );
  NOR2_X1 U12 ( .A1(d__apx[11]), .A2(acc__sel), .ZN(n12) );
  AOI21_X1 U13 ( .B1(d__acc[27]), .B2(acc__sel), .A(n12), .ZN(\d[27]_BAR ) );
  NOR2_X1 U14 ( .A1(n5), .A2(acc__sel), .ZN(n14) );
  AOI21_X1 U15 ( .B1(d__acc[28]), .B2(acc__sel), .A(n14), .ZN(\d[28]_BAR ) );
  NAND2_X1 U16 ( .A1(d__acc[29]), .A2(acc__sel), .ZN(n16) );
  OAI21_X1 U17 ( .B1(d__apx[13]), .B2(acc__sel), .A(n16), .ZN(d[29]) );
  NAND2_X1 U18 ( .A1(d__acc[30]), .A2(acc__sel), .ZN(n17) );
  OAI21_X1 U19 ( .B1(d__apx[14]), .B2(acc__sel), .A(n17), .ZN(d[30]) );
  NAND2_X1 U20 ( .A1(d__acc[31]), .A2(acc__sel), .ZN(n18) );
  OAI21_X1 U21 ( .B1(d__apx[15]), .B2(acc__sel), .A(n18), .ZN(d[31]) );
  MUX2_X1 U22 ( .A(d__apx[16]), .B(d__acc[32]), .S(acc__sel), .Z(d[32]) );
  NAND2_X1 U23 ( .A1(d__acc[33]), .A2(acc__sel), .ZN(n19) );
  OAI21_X1 U24 ( .B1(d__apx[17]), .B2(acc__sel), .A(n19), .ZN(d[33]) );
  MUX2_X1 U25 ( .A(d__apx[18]), .B(d__acc[34]), .S(acc__sel), .Z(d[34]) );
  MUX2_X1 U26 ( .A(d__apx[19]), .B(d__acc[35]), .S(acc__sel), .Z(d[35]) );
  MUX2_X1 U27 ( .A(d__apx[20]), .B(d__acc[36]), .S(acc__sel), .Z(d[36]) );
  MUX2_X1 U28 ( .A(d__apx[21]), .B(d__acc[37]), .S(acc__sel), .Z(d[37]) );
  NAND2_X1 U29 ( .A1(d__acc[38]), .A2(acc__sel), .ZN(n20) );
  OAI21_X1 U30 ( .B1(d__apx[22]), .B2(acc__sel), .A(n20), .ZN(d[38]) );
  NAND2_X1 U31 ( .A1(d__acc[39]), .A2(acc__sel), .ZN(n21) );
  OAI21_X1 U32 ( .B1(d__apx[23]), .B2(acc__sel), .A(n21), .ZN(d[39]) );
  NAND2_X1 U33 ( .A1(d__acc[40]), .A2(acc__sel), .ZN(n22) );
  OAI21_X1 U34 ( .B1(d__apx[24]), .B2(acc__sel), .A(n22), .ZN(d[40]) );
  MUX2_X1 U35 ( .A(d__apx[25]), .B(d__acc[41]), .S(acc__sel), .Z(d[41]) );
  NAND2_X1 U36 ( .A1(d__acc[42]), .A2(acc__sel), .ZN(n23) );
  OAI21_X1 U37 ( .B1(d__apx[26]), .B2(acc__sel), .A(n23), .ZN(d[42]) );
  NAND2_X1 U38 ( .A1(d__acc[43]), .A2(acc__sel), .ZN(n24) );
  OAI21_X1 U39 ( .B1(d__apx[27]), .B2(acc__sel), .A(n24), .ZN(d[43]) );
  MUX2_X1 U40 ( .A(d__apx[28]), .B(d__acc[44]), .S(acc__sel), .Z(d[44]) );
  MUX2_X1 U41 ( .A(d__apx[29]), .B(d__acc[45]), .S(acc__sel), .Z(d[45]) );
  MUX2_X1 U42 ( .A(d__apx[30]), .B(d__acc[46]), .S(acc__sel), .Z(d[46]) );
  MUX2_X1 U43 ( .A(d__apx[31]), .B(d__acc[47]), .S(acc__sel), .Z(d[47]) );
  MUX2_X1 U44 ( .A(d__apx[32]), .B(d__acc[48]), .S(acc__sel), .Z(d[48]) );
  NAND2_X1 U45 ( .A1(d__acc[49]), .A2(acc__sel), .ZN(n25) );
  OAI21_X1 U46 ( .B1(d__apx[33]), .B2(acc__sel), .A(n25), .ZN(d[49]) );
  MUX2_X1 U47 ( .A(d__apx[34]), .B(d__acc[50]), .S(acc__sel), .Z(d[50]) );
  MUX2_X1 U48 ( .A(d__apx[35]), .B(d__acc[51]), .S(acc__sel), .Z(d[51]) );
  NAND2_X1 U49 ( .A1(d__acc[52]), .A2(acc__sel), .ZN(n26) );
  OAI21_X1 U50 ( .B1(d__apx[36]), .B2(acc__sel), .A(n26), .ZN(d[52]) );
  NAND2_X1 U51 ( .A1(d__acc[53]), .A2(acc__sel), .ZN(n27) );
  OAI21_X1 U52 ( .B1(d__apx[37]), .B2(acc__sel), .A(n27), .ZN(d[53]) );
  NAND2_X1 U53 ( .A1(d__acc[54]), .A2(acc__sel), .ZN(n28) );
  OAI21_X1 U54 ( .B1(d__apx[38]), .B2(acc__sel), .A(n28), .ZN(d[54]) );
  NAND2_X1 U55 ( .A1(d__acc[55]), .A2(acc__sel), .ZN(n29) );
  OAI21_X1 U56 ( .B1(d__apx[39]), .B2(acc__sel), .A(n29), .ZN(d[55]) );
  MUX2_X1 U57 ( .A(d__apx[40]), .B(d__acc[56]), .S(acc__sel), .Z(d[56]) );
  NAND2_X1 U58 ( .A1(d__acc[57]), .A2(acc__sel), .ZN(n30) );
  OAI21_X1 U59 ( .B1(d__apx[41]), .B2(acc__sel), .A(n30), .ZN(d[57]) );
  NAND2_X1 U60 ( .A1(d__acc[58]), .A2(acc__sel), .ZN(n31) );
  OAI21_X1 U61 ( .B1(d__apx[42]), .B2(acc__sel), .A(n31), .ZN(d[58]) );
  MUX2_X1 U62 ( .A(d__apx[43]), .B(d__acc[59]), .S(acc__sel), .Z(d[59]) );
  MUX2_X1 U63 ( .A(d__apx[44]), .B(d__acc[60]), .S(acc__sel), .Z(d[60]) );
  NAND2_X1 U64 ( .A1(d__acc[61]), .A2(acc__sel), .ZN(n32) );
  OAI21_X1 U65 ( .B1(d__apx[45]), .B2(acc__sel), .A(n32), .ZN(d[61]) );
  NAND2_X1 U66 ( .A1(d__acc[62]), .A2(acc__sel), .ZN(n33) );
  OAI21_X1 U67 ( .B1(d__apx[46]), .B2(acc__sel), .A(n33), .ZN(d[62]) );
  MUX2_X1 U68 ( .A(d__apx[47]), .B(d__acc[63]), .S(acc__sel), .Z(d[63]) );
  NAND2_X1 U69 ( .A1(acc__sel), .A2(d__acc[21]), .ZN(n34) );
  OAI21_X1 U70 ( .B1(d__apx[5]), .B2(acc__sel), .A(n34), .ZN(d[21]) );
  NAND2_X1 U71 ( .A1(acc__sel), .A2(d__acc[22]), .ZN(n35) );
  OAI21_X1 U72 ( .B1(n3), .B2(acc__sel), .A(n35), .ZN(d[22]) );
  NAND2_X1 U73 ( .A1(acc__sel), .A2(d__acc[23]), .ZN(n36) );
  OAI21_X1 U74 ( .B1(n4), .B2(acc__sel), .A(n36), .ZN(d[23]) );
  NAND2_X1 U75 ( .A1(acc__sel), .A2(d__acc[20]), .ZN(n37) );
  OAI21_X1 U76 ( .B1(d__apx[4]), .B2(acc__sel), .A(n37), .ZN(d[20]) );
  AND2_X1 U77 ( .A1(acc__sel), .A2(d__acc[0]), .ZN(d[0]) );
  AND2_X1 U78 ( .A1(acc__sel), .A2(d__acc[1]), .ZN(d[1]) );
  AND2_X1 U79 ( .A1(acc__sel), .A2(d__acc[2]), .ZN(d[2]) );
  AND2_X1 U80 ( .A1(acc__sel), .A2(d__acc[3]), .ZN(d[3]) );
  AND2_X1 U81 ( .A1(acc__sel), .A2(d__acc[4]), .ZN(d[4]) );
  AND2_X1 U82 ( .A1(acc__sel), .A2(d__acc[5]), .ZN(d[5]) );
  AND2_X1 U83 ( .A1(acc__sel), .A2(d__acc[6]), .ZN(d[6]) );
  AND2_X1 U84 ( .A1(acc__sel), .A2(d__acc[7]), .ZN(d[7]) );
  AND2_X1 U85 ( .A1(acc__sel), .A2(d__acc[8]), .ZN(d[8]) );
  AND2_X1 U86 ( .A1(acc__sel), .A2(d__acc[9]), .ZN(d[9]) );
  AND2_X1 U87 ( .A1(acc__sel), .A2(d__acc[10]), .ZN(d[10]) );
  AND2_X1 U88 ( .A1(acc__sel), .A2(d__acc[11]), .ZN(d[11]) );
  AND2_X1 U89 ( .A1(acc__sel), .A2(d__acc[12]), .ZN(d[12]) );
  AND2_X1 U90 ( .A1(acc__sel), .A2(d__acc[13]), .ZN(d[13]) );
  AND2_X1 U91 ( .A1(acc__sel), .A2(d__acc[14]), .ZN(d[14]) );
  AND2_X1 U92 ( .A1(acc__sel), .A2(d__acc[15]), .ZN(d[15]) );
  MUX2_X1 U93 ( .A(d__apx[0]), .B(d__acc[16]), .S(acc__sel), .Z(d[16]) );
  MUX2_X1 U94 ( .A(d__apx[1]), .B(d__acc[17]), .S(acc__sel), .Z(d[17]) );
  MUX2_X1 U95 ( .A(d__apx[2]), .B(d__acc[18]), .S(acc__sel), .Z(d[18]) );
  MUX2_X1 U96 ( .A(n2), .B(d__acc[19]), .S(acc__sel), .Z(\d[19] ) );
  conf_int_mul__noFF__arch_agnos_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 mul__inst ( 
        .clk(clk), .rst(n1), .a(a), .b(b), .\d[47] (d__apx[47]), .\d[44] (
        d__apx[44]), .\d[43] (d__apx[43]), .\d[40] (d__apx[40]), .\d[37]_BAR (
        d__apx[37]), .\d[34] (d__apx[34]), .\d[31] (d__apx[31]), .\d[28] (
        d__apx[28]), .\d[16] (d__apx[16]), .\d[1] (d__apx[1]), .\d[0] (
        d__apx[0]), .\d[33]_BAR (d__apx[33]), .\d[27]_BAR (d__apx[27]), 
        .\d[26]_BAR (d__apx[26]), .\d[24]_BAR (d__apx[24]), .\d[23]_BAR (
        d__apx[23]), .\d[15]_BAR (d__apx[15]), .\d[14]_BAR (d__apx[14]), 
        .\d[11]_BAR (d__apx[11]), .\d[9]_BAR (d__apx[9]), .\d[4]_BAR (
        d__apx[4]), .\d[42]_BAR (d__apx[42]), .\d[41]_BAR (d__apx[41]), 
        .\d[30] (d__apx[30]), .\d[22]_BAR (d__apx[22]), .\d[46]_BAR (
        d__apx[46]), .\d[35] (d__apx[35]), .\d[19] (d__apx[19]), .\d[10]_BAR (
        d__apx[10]), .\d[8]_BAR (d__apx[8]), .\d[5]_BAR (d__apx[5]), .\d[29] (
        d__apx[29]), .\d[32] (d__apx[32]), .\d[39]_BAR (d__apx[39]), .\d[2] (
        d__apx[2]), .\d[36]_BAR (d__apx[36]), .\d[25] (d__apx[25]), 
        .\d[13]_BAR (d__apx[13]), .\d[38]_BAR (d__apx[38]), .\d[20] (
        d__apx[20]), .\d[18] (d__apx[18]), .\d[17]_BAR (d__apx[17]), 
        .\d[45]_BAR (d__apx[45]), .\d[21] (d__apx[21]), .\d[12] (d__apx[12]), 
        .\d[7] (d__apx[7]), .\d[6] (d__apx[6]), .\d[3]_BAR (d__apx[3]) );
endmodule
