library verilog;
use verilog.vl_types.all;
entity UDP_typical_MGM_H_IQ_FF_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end UDP_typical_MGM_H_IQ_FF_UDP;
