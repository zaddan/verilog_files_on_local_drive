library verilog;
use verilog.vl_types.all;
entity OAI221_X1_func is
    port(
        A               : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        C1              : in     vl_logic;
        C2              : in     vl_logic;
        ZN              : out    vl_logic
    );
end OAI221_X1_func;
