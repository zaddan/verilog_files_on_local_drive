module conf_int_mul__noFF__arch_agnos_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 ( clk, 
        rst, a, b, \d[47] , \d[44] , \d[43] , \d[40] , \d[37]_BAR , \d[34] , 
        \d[31] , \d[28] , \d[16] , \d[1] , \d[0] , \d[33]_BAR , \d[27]_BAR , 
        \d[26]_BAR , \d[24]_BAR , \d[23]_BAR , \d[21]_BAR , \d[15]_BAR , 
        \d[14]_BAR , \d[11]_BAR , \d[9]_BAR , \d[6]_BAR , \d[4]_BAR , 
        \d[42]_BAR , \d[41]_BAR , \d[30] , \d[22]_BAR , \d[46]_BAR , \d[35] , 
        \d[19] , \d[10]_BAR , \d[8]_BAR , \d[5]_BAR , \d[3] , \d[29] , 
        \d[7]_BAR , \d[32] , \d[39]_BAR , \d[12]_BAR , \d[2] , \d[36]_BAR , 
        \d[25] , \d[13]_BAR , \d[38]_BAR , \d[20] , \d[18] , \d[45] , 
        \d[17]_BAR  );
  input [23:0] a;
  input [23:0] b;
  input clk, rst;
  output \d[47] , \d[44] , \d[43] , \d[40] , \d[37]_BAR , \d[34] , \d[31] ,
         \d[28] , \d[16] , \d[1] , \d[0] , \d[33]_BAR , \d[27]_BAR ,
         \d[26]_BAR , \d[24]_BAR , \d[23]_BAR , \d[21]_BAR , \d[15]_BAR ,
         \d[14]_BAR , \d[11]_BAR , \d[9]_BAR , \d[6]_BAR , \d[4]_BAR ,
         \d[42]_BAR , \d[41]_BAR , \d[30] , \d[22]_BAR , \d[46]_BAR , \d[35] ,
         \d[19] , \d[10]_BAR , \d[8]_BAR , \d[5]_BAR , \d[3] , \d[29] ,
         \d[7]_BAR , \d[32] , \d[39]_BAR , \d[12]_BAR , \d[2] , \d[36]_BAR ,
         \d[25] , \d[13]_BAR , \d[38]_BAR , \d[20] , \d[18] , \d[45] ,
         \d[17]_BAR ;
  wire   n5798, n976, n5808, n5807, n5838, n2157, n5918, n4973, n5610, n5609,
         n369, n1243, n989, n4583, n1634, n5036, n5091, n1756, n1755, n3125,
         n690, n3409, n520, n521, n4907, n4281, n4282, n2114, n3158, n5357,
         n5556, n1150, n1152, n5694, n3245, n3248, n4906, n604, n605, n3561,
         n3421, n3824, n3823, n2170, n2523, n3023, n1863, n1862, n2201, n811,
         n812, n557, n5359, n5358, n5457, n3237, n3475, n3747, n5079, n3540,
         n1225, n2871, n2874, n2870, n3251, n4741, n2314, n2103, n4743, n1960,
         n1193, n3217, n1397, n1646, n1647, n2076, n463, n464, n2836, n461,
         n2828, n3915, n3916, n159, n1477, n3404, n4692, n4762, n5075, n947,
         n3242, n3241, n5167, n4239, n4217, n4788, n2596, n1287, n4100, n923,
         n3435, n1554, n921, n5294, n5190, n3760, n4607, n865, n3533, n3642,
         n4770, n3617, n3324, n2717, n3562, n2270, n1147, n4489, n3757, n3209,
         n5477, n5947, n984, n4677, n1064, n29, n1194, n635, n981, n513, n1329,
         n734, n3952, n4733, n753, n3220, n1847, n5293, n2412, n194, n911,
         n5718, n2305, n304, n614, n5413, n5412, n5541, n5414, n2043, n4952,
         n808, n2093, n949, n1633, n5514, n5513, n5547, n5235, n2914, n2744,
         n2715, n4834, n5074, n5951, n2116, n2309, n2786, n2933, n5376, n2785,
         n5119, n5117, n5197, n1981, n3369, n529, n528, n6093, n2700, n4777,
         n2256, n3882, n3881, n3883, n328, n4559, n1, n2, n394, n1411, n392,
         n5300, n3, n3985, n3813, n3814, n4, n391, n1406, n5184, n564, n5185,
         n5242, n5241, n5240, n5303, n5169, n5, n6, n5168, n1999, n1429, n1430,
         n283, n1534, n2189, n3149, n4480, n7, n8, n1093, n170, n2184, n4463,
         n1852, n2548, n3755, n1851, n1408, n971, n1407, n5308, n1019, n2430,
         n2274, n2275, n2137, n4051, n4118, n4490, n6183, n4142, n3856, n3855,
         n3898, n3730, n4333, n4332, n2124, n11, n4450, n3042, n14, n13, n6149,
         n4472, n3265, n909, n4527, n251, n3957, n4034, n3894, n1050, n1432,
         n261, n262, n264, n3049, n3050, n15, n4363, n2009, n16, n174, n941,
         n1583, n2909, n2910, n2912, n6336, n5834, n2006, n5323, n1051, n2104,
         n3802, n17, n3694, n3693, n3307, n2187, n1363, n1362, n1973, n4496,
         n2511, n2868, n2869, n4478, n3446, n2566, n4085, n813, n816, n4350,
         n4351, n4349, n3308, n4354, n21, n20, n3072, n4405, n2411, n674, n22,
         n323, n3234, n321, n4566, n4267, n4266, n5699, n23, n288, n4254,
         n1582, n1581, n4557, n24, n27, n25, n5776, n5774, n6454, n771, n5725,
         n2031, n4565, n760, n4734, n30, n1571, n3283, n651, n2283, n3468,
         n1470, n4319, n4318, n2676, n1008, n6187, n1117, n2229, n31, n4636,
         n2375, n6366, n3069, n3070, n4040, n3197, n3196, n1831, n869, n868,
         n5629, n2003, n584, n1469, n3753, n3645, n2215, n1700, n866, n1702,
         n1701, n4465, n32, n444, n1333, n442, n443, n1483, n1482, n633, n5252,
         n2291, n871, n4061, n4055, n4057, n4601, n3606, n5188, n1394, n1390,
         n5239, n1391, n5151, n4781, n33, n4785, n5260, n454, n37, n5174,
         n5173, n1042, n38, n2518, n1088, n2826, n2410, n6214, n1041, n5930,
         n259, n6134, n5255, n5253, n5171, n5172, n39, n5295, n41, n6513,
         n4895, n433, n1060, n805, n2143, n1980, n1107, n4614, n1191, n44,
         n661, n2398, n659, n660, n4824, n1063, n2371, n45, n5555, n1724,
         n5557, n2520, n2522, n5094, n3466, n2767, n6221, n2644, n49, n2692,
         n2694, n2769, n562, n561, n1996, n4650, n1994, n2693, n1846, n3126,
         n5804, n3672, n1079, n1667, n3602, n3603, n1081, n1080, n50, n5320,
         n5596, n5919, n628, n343, n1985, n1984, n4912, n895, n894, n337,
         n4071, n1295, n1294, n4759, n4758, n2321, n1788, n3869, n4219, n3912,
         n3448, n3447, n2374, n51, n3482, n2110, n2111, n485, n3706, n3745,
         n1458, n3521, n3523, n3350, n1641, n3524, n53, n6151, n1338, n3491,
         n281, n2298, n3983, n2238, n3304, n54, n55, n3289, n2383, n697, n696,
         n2473, n6000, n5616, n6200, n1943, n172, n4882, n1440, n2583, n3474,
         n3396, n699, n3538, n1933, n4073, n819, n2500, n2849, n3557, n3011,
         n5360, n2502, n6654, n245, n993, n4890, n59, n4921, n4889, n1798,
         n1800, n5019, n824, n823, n1507, n2757, n60, n6086, n61, n3161, n3342,
         n1102, n2326, n4558, n1276, n1775, n1774, n1773, n4657, n2546, n3130,
         n3129, n3127, n6450, n1457, n4529, n4408, n2995, n4042, n63, n3775,
         n3776, n66, n3778, n6161, n6445, n1911, n1910, n1913, n1912, n3654,
         n69, n2508, n4231, n70, n71, n4338, n2180, n4488, n990, n2081, n72,
         n1140, n6186, n2602, n73, n349, n4069, n347, n348, n3052, n4582,
         n2130, n2167, n74, n4300, n4298, n1320, n5717, n4296, n4297, n75,
         n1914, n78, n779, n3073, n777, n4721, n4578, n4577, n4580, n1759,
         n5212, n4514, n4517, n758, n2249, n3175, n1448, n4356, n80, n4404,
         n83, n81, n4598, n5471, n5364, n3285, n1976, n3078, n84, n2235, n86,
         n1753, n1754, n4479, n4584, n1997, n3650, n3901, n2649, n4637, n4635,
         n2226, n1110, n4476, n998, n87, n757, n756, n3064, n88, n2090, n1157,
         n3731, n2131, n2092, n2324, n754, n279, n278, n89, n4005, n4293,
         n3941, n6558, n91, n4056, n94, n92, n4506, n95, n791, n793, n3974,
         n992, n988, n3904, n4376, n2347, n432, n2929, n931, n4515, n4512,
         n2325, n4612, n3568, n96, n1848, n2469, n1417, n525, n524, n1077, n98,
         n2243, n319, n930, n101, n100, n2818, n2491, n254, n4670, n2156,
         n1098, n2152, n1710, n2042, n3331, n2646, n4563, n4564, n1006, n3408,
         n2803, n1004, n4486, n3051, n4576, n6402, n676, n677, n5324, n103,
         n5027, n6452, n2750, n1619, n1035, n6022, n1145, n6023, n1781, n1780,
         n5111, n1779, n6569, n3664, n1506, n5210, n509, n2749, n3624, n4689,
         n4816, n4924, n611, n585, n2272, n108, n5032, n5038, n2600, n2599,
         n1540, n1685, n875, n2063, n1721, n2064, n2810, n5929, n2330, n5926,
         n6005, n1675, n916, n1024, n2218, n809, n810, n111, n110, n1907,
         n1941, n5039, n1112, n1942, n4604, n3085, n4481, n1127, n1930, n116,
         n114, n113, n2406, n1992, n1991, n117, n1380, n1336, n418, n419,
         n5277, n118, n737, n738, n119, n3500, n646, n120, n787, n2530, n2331,
         n388, n123, n4528, n1600, n2691, n2690, n3832, n2276, n1957, n124,
         n4838, n1224, n4839, n1226, n2348, n2051, n2050, n125, n1270, n127,
         n3670, n5862, n2879, n5867, n5314, n3105, n2044, n5069, n2468, n1285,
         n132, n2295, n3937, n3938, n280, n2517, n5133, n133, n5014, n136,
         n134, n5058, n6035, n137, n691, n1716, n689, n1714, n1530, n6391,
         n1713, n1240, n4901, n2219, n595, n594, n256, n6525, n3758, n5593,
         n4805, n139, n2936, n5389, n5388, n1164, n1163, n4760, n1091, n141,
         n140, n3275, n142, n1321, n1925, n5729, n143, n1752, n1594, n4589,
         n1529, n2470, n3727, n4720, n1437, n4656, n4655, n1339, n5886, n145,
         n6062, n5876, n5884, n4736, n146, n1350, n1376, n4975, n2949, n5839,
         n2975, n2974, n4917, n573, n1375, n2488, n1653, n3253, n3713, n148,
         n2384, n1844, n150, n149, n1845, n1683, n4904, n4905, n3074, n3077,
         n6202, n3273, n1461, n5099, n5377, n154, n2630, n3247, n3080, n4539,
         n6377, n2852, n1947, n3157, n6059, n6055, n3726, n2278, n4599, n586,
         n1546, n1202, n162, n1850, n1465, n5647, n163, n3113, n3114, n1500,
         n1502, n1501, n217, n4592, n2313, n2315, n4833, n3385, n3469, n2643,
         n2642, n164, n165, n5392, n5393, n5391, n1327, n345, n5390, n3724,
         n3359, n4982, n4409, n4410, n4411, n4412, n4070, n818, n2973, n2510,
         n2382, n5034, n166, n2597, n3090, n3089, n5458, n1344, n167, n5995,
         n6068, n5931, n5508, n972, n2069, n169, n168, n5553, n5552, n1267,
         n1265, n3155, n1778, n952, n538, n780, n214, n2403, n1769, n4651,
         n4735, n4520, n4519, n4573, n192, n1504, n1176, n173, n3986, n1175,
         n3984, n4277, n4279, n2208, n3843, n3842, n3009, n1257, n3008, n1149,
         n2506, n939, n940, n3076, n6587, n2847, n1013, n5984, n5973, n657,
         n658, n4158, n175, n4247, n4285, n1551, n1553, n4245, n2172, n268,
         n620, n619, n5305, n176, n5302, n5301, n3286, n4295, n2831, n2669,
         n2668, n2964, n2963, n177, n339, n178, n387, n386, n548, n179, n550,
         n2971, n1136, n1355, n5975, n5970, n2099, n3024, n448, n5143, n5056,
         n181, n4194, n4193, n4192, n5689, n183, n182, n5139, n5136, n2248,
         n1969, n1038, n3211, n857, n3591, n4307, n2242, n2241, n3364, n2173,
         n842, n4229, n4228, n1123, n3588, n3589, n2388, n3213, n2389, n1200,
         n1197, n4667, n1279, n1280, n2179, n190, n4470, n2366, n3853, n3852,
         n3892, n1159, n1158, n3303, n195, n1873, n1370, n601, n3095, n3087,
         n4469, n1842, n196, n731, n3192, n729, n5558, n5924, n3389, n4977,
         n197, n2458, n2457, n2460, n2467, n3457, n4183, n3456, n199, n198,
         n4185, n202, n201, n4353, n4346, n1603, n5894, n5554, n5562, n4995,
         n6158, n4401, n1932, n4794, n4810, n206, n5055, n1515, n1516, n1517,
         n282, n5053, n1749, n1748, n1747, n1639, n1638, n5049, n5047, n5045,
         n5042, n5044, n510, n1627, n327, n208, n1962, n4075, n1961, n3980,
         n2972, n6017, n5381, n6205, n6021, n979, n1974, n2421, n3877, n3975,
         n792, n978, n3636, n3635, n5144, n2108, n3991, n211, n210, n2005,
         n788, n789, n4484, n1468, n1467, n664, n213, n702, n4776, n700, n701,
         n892, n4869, n2182, n2181, n215, n1027, n2163, n2083, n3580, n2117,
         n3264, n216, n1511, n2166, n2479, n2601, n3086, n4545, n4624, n218,
         n655, n653, n654, n1612, n5489, n1610, n2540, n5451, n5450, n5452,
         n5506, n1179, n221, n219, n5276, n309, n223, n222, n5342, n4767, n566,
         n2435, n2434, n2524, n2032, n3263, n3481, n2926, n2917, n2426, n1599,
         n4908, n4909, n5369, n2812, n2072, n5546, n621, n622, n228, n652,
         n3083, n4365, n4012, n229, n1988, n4740, n4821, n4668, n232, n3221,
         n2969, n3407, n3551, n3388, n1274, n3552, n3553, n3872, n253, n3871,
         n3911, n234, n1833, n1832, n1835, n1834, n235, n2461, n1665, n1022,
         n2837, n1266, n236, n852, n5764, n850, n851, n4474, n534, n3417,
         n3418, n3420, n238, n1185, n6446, n3571, n265, n239, n6614, n5326,
         n1016, n2086, n4641, n4640, n243, n241, n5361, n4829, n5526, n1212,
         n5076, n4502, n745, n744, n244, n5566, n5564, n1723, n3215, n4550,
         n1882, n4674, n4130, n246, n4135, n249, n247, n4216, n248, n1009,
         n2952, n4316, n260, n5322, n1324, n2526, n3208, n255, n4549, n5105,
         n4526, n257, n827, n828, n258, n1909, n4315, n2334, n2721, n263,
         n2707, n4007, n712, n2223, n4375, n4837, n2834, n2956, n4686, n1509,
         n3900, n266, n3903, n3554, n270, n272, n662, n663, n665, n6206, n4972,
         n274, n1343, n2107, n275, n276, n430, n2337, n5996, n6070, n4551,
         n4552, n4669, n2513, n4754, n5010, n3656, n3705, n3453, n4212, n4746,
         n4214, n2770, n2550, n4248, n1865, n4001, n3811, n3809, n3555, n1964,
         n4077, n1963, n1412, n2783, n2784, n2779, n1868, n5789, n290, n4605,
         n1218, n4608, n3860, n3861, n4913, n2731, n4322, n4323, n293, n3756,
         n6160, n2333, n297, n298, n296, n300, n301, n303, n3075, n1181, n6029,
         n5895, n4437, n3942, n2587, n307, n305, n306, n308, n3976, n4939,
         n1479, n4314, n1431, n311, n2743, n1565, n4447, n317, n318, n4466,
         n1075, n3959, n3958, n3961, n3683, n4899, n2987, n2373, n320, n4009,
         n4998, n4392, n4394, n2738, n3700, n3945, n2300, n324, n3235, n1826,
         n1825, n326, n2391, n1082, n4131, n4188, n4189, n5070, n5287, n5355,
         n331, n329, n330, n332, n5331, n3704, n4704, n1790, n3581, n3600,
         n4919, n3575, n2752, n4979, n4976, n5851, n4780, n3313, n4779, n4962,
         n3886, n5149, n2358, n2357, n2489, n2355, n333, n334, n336, n4038,
         n4504, n3329, n4499, n4498, n3430, n338, n3190, n3870, n1012, n1735,
         n4933, n4811, n5307, n5317, n340, n2251, n2254, n341, n4370, n3695,
         n342, n881, n1609, n5572, n5913, n1099, n5384, n1776, n4457, n4019,
         n351, n4289, n4288, n4287, n4302, n4903, n354, n360, n466, n359, n361,
         n1720, n1719, n365, n672, n673, n366, n1000, n367, n3154, n1261,
         n1260, n368, n5888, n1715, n372, n370, n371, n373, n2629, n2066, n376,
         n374, n375, n377, n4871, n2651, n4452, n380, n378, n4025, n1874,
         n3338, n3337, n4628, n3336, n2537, n383, n3438, n5266, n384, n5459,
         n385, n2329, n5298, n5297, n395, n4703, n4994, n4434, n4989, n2809,
         n489, n3917, n4568, n4569, n5084, n1830, n2594, n5024, n985, n3088,
         n2397, n5176, n2401, n1629, n1765, n397, n3981, n3982, n3923, n2843,
         n3323, n4769, n400, n401, n4407, n4406, n4413, n3919, n4059, n405,
         n3943, n4065, n406, n3166, n2010, n2322, n3939, n1746, n5155, n409,
         n407, n408, n410, n3403, n412, n413, n5072, n414, n1455, n4058, n4064,
         n3944, n1259, n1258, n1148, n415, n1484, n4524, n416, n2102, n3492,
         n4914, n2613, n5672, n3722, n421, n5667, n422, n4099, n424, n425,
         n434, n4845, n5952, n4812, n4814, n581, n830, n832, n4856, n4863,
         n1556, n3461, n5707, n3362, n4050, n4442, n6015, n6014, n3476, n6019,
         n2230, n2231, n1545, n4942, n3994, n5620, n6016, n2724, n470, n4775,
         n3204, n2038, n435, n493, n716, n437, n438, n468, n441, n817, n3831,
         n650, n4966, n5092, n2928, n3370, n2853, n6596, n1071, n1023, n5332,
         n5334, n446, n1596, n1595, n452, n3108, n1379, n3817, n3816, n3820,
         n3815, n2151, n2153, n4974, n821, n822, n458, n3570, n5875, n5868,
         n4874, n459, n4630, n4866, n2639, n460, n3867, n1436, n1387, n4389,
         n531, n5840, n1510, n5611, n5453, n5999, n1607, n5491, n5490, n5493,
         n755, n2889, n4342, n3736, n2563, n471, n472, n2054, n2811, n5368,
         n6504, n3355, n4309, n2927, n2918, n3792, n2199, n2198, n3887, n4774,
         n3935, n3936, n3934, n588, n4654, n591, n2758, n2516, n2515, n2830,
         n2603, n2310, n1544, n1543, n477, n4372, n480, n478, n479, n481,
         n5449, n482, n2303, n483, n484, n6031, n6030, n6028, n6122, n4473,
         n5035, n556, n2925, n5529, n2923, n5916, n5678, n3153, n3188, n647,
         n1263, n486, n2196, n490, n488, n491, n3586, n747, n761, n750, n3545,
         n522, n4920, n494, n492, n5059, n831, n3160, n499, n498, n503, n504,
         n1978, n501, n502, n4078, n4080, n4865, n4864, n2640, n505, n506,
         n507, n508, n815, n511, n5220, n3504, n3684, n512, n515, n514, n517,
         n518, n519, n4867, n523, n4763, n530, n2267, n2268, n710, n2155,
         n5828, n2200, n1299, n267, n1886, n1768, n4475, n536, n537, n2638,
         n6325, n2637, n1435, n1434, n5341, n1153, n1154, n539, n2865, n1927,
         n3465, n2746, n2161, n1920, n3239, n3063, n4581, n5621, n1840, n5792,
         n3367, n1687, n2339, n542, n540, n541, n4205, n546, n544, n1137, n549,
         n5676, n2519, n102, n553, n551, n552, n554, n5031, n563, n6607, n4642,
         n2039, n5040, n3431, n975, n559, n560, n4662, n2967, n4661, n2695,
         n1059, n4586, n1083, n1628, n571, n572, n4916, n575, n574, n576,
         n2327, n4997, n3631, n2512, n4046, n3620, n2902, n2129, n648, n2128,
         n1360, n1549, n3996, n1550, n1871, n4795, n606, n4211, n2101, n2699,
         n2968, n6204, n593, n4802, n598, n599, n3150, n2336, n4606, n600,
         n2082, n602, n603, n6207, n1870, n3315, n5817, n2154, n1104, n5023,
         n3305, n4348, n608, n4554, n4555, n2806, n1881, n609, n2253, n3450,
         n3622, n2354, n1875, n1813, n1805, n1812, n4570, n4232, n3296, n5374,
         n3663, n5853, n4483, n2950, n1151, n5660, n4150, n4149, n688, n2932,
         n615, n3746, n6331, n5383, n616, n1031, n1505, n1120, n2438, n617,
         n618, n5275, n5345, n465, n3691, n4633, n4632, n4631, n1076, n6610,
         n4402, n4523, n5112, n999, n1622, n1674, n626, n627, n5472, n624,
         n625, n5525, n1709, n951, n436, n1660, n629, n4959, n749, n5991,
         n5983, n5982, n5989, n4373, n3738, n4969, n630, n5218, n4320, n4731,
         n4730, n934, n933, n5217, n5206, n5216, n637, n5630, n5120, n5118,
         n5177, n2538, n2539, n642, n640, n641, n643, n5780, n3833, n3029,
         n5077, n5336, n1745, n1744, n2195, n2437, n766, n4072, n3913, n6527,
         n943, n4511, n4510, n2788, n3201, n2913, n1946, n995, n3318, n5897,
         n3351, n2096, n6529, n1880, n3954, n3368, n3953, n3955, n3202, n3082,
         n4382, n2296, n3015, n314, n1190, n5427, n5437, n1598, n649, n2824,
         n4671, n1105, n1698, n5330, n1785, n668, n675, n1002, n3625, n4753,
         n4752, n3278, n4308, n4244, n678, n679, n1741, n1351, n5870, n682,
         n683, n681, n5043, n687, n686, n3530, n5869, n4968, n1215, n1230,
         n3259, n3258, n705, n706, n5041, n703, n3587, n1937, n4684, n707,
         n2578, n2588, n5745, n5768, n5769, n1898, n3680, n1986, n1134, n1133,
         n3452, n4037, n3594, n2368, n3060, n2367, n4961, n714, n4964, n713,
         n715, n2576, n6511, n2883, n4339, n6609, n5288, n5289, n719, n6152,
         n6150, n720, n5238, n1877, n723, n721, n722, n724, n4999, n3056,
         n1564, n5424, n6515, n3020, n2408, n3907, n3191, n727, n725, n5563,
         n728, n1284, n1066, n733, n735, n3573, n1524, n5315, n3371, n736,
         n2930, n4575, n739, n3838, n3764, n4271, n3462, n3834, n3266, n2846,
         n5354, n742, n740, n741, n743, n2813, n746, n473, n2899, n1694, n4067,
         n748, n3509, n3346, n751, n1281, n3836, n4335, n2146, n2589, n2954,
         n5670, n5671, n5677, n1993, n2719, n1727, n4854, n4862, n4855, n1378,
         n759, n937, n833, n4705, n2658, n2882, n3930, n3932, n764, n763,
         n1593, n769, n767, n3896, n3895, n967, n1010, n772, n773, n775, n2087,
         n4649, n4737, n2311, n2773, n4538, n807, n781, n4159, n2097, n4161,
         n2246, n2245, n782, n1039, n3928, n2444, n2074, n2073, n785, n784,
         n1983, n3528, n3529, n790, n3522, n1637, n1836, n1201, n3607, n3598,
         n3284, n2839, n3013, n800, n802, n4652, n803, n804, n3480, n4435,
         n2159, n4900, n1300, n5090, n5089, n2799, n4145, n4144, n4143, n5658,
         n3224, n964, n1113, n2562, n2559, n2561, n5665, n4152, n4151, n3905,
         n2307, n6456, n3131, n1322, n825, n826, n6514, n980, n5060, n2544,
         n4000, n838, n836, n837, n839, n845, n843, n844, n846, n3395, n4387,
         n4388, n1141, n4175, n1626, n4197, n1783, n2360, n1782, n5113, n5777,
         n5765, n5772, n2113, n855, n853, n854, n856, n3325, n1630, n4724,
         n860, n2239, n4275, n863, n861, n862, n6608, n4796, n3463, n2140,
         n4272, n3806, n6215, n3807, n867, n870, n873, n877, n880, n3219,
         n3291, n3290, n3268, n1858, n1903, n1905, n3854, n2748, n2168, n1247,
         n2683, n2682, n4765, n6519, n882, n2966, n885, n2205, n5246, n889,
         n887, n3868, n2308, n891, n1223, n2084, n2085, n6655, n2543, n3365,
         n903, n1124, n2077, n2369, n4872, n914, n912, n913, n915, n1025, n919,
         n917, n918, n920, n5883, n925, n926, n928, n927, n2004, n932, n5571,
         n5373, n2323, n2720, n4509, n1935, n944, n4593, n4726, n4681, n4749,
         n4611, n3292, n4880, n1864, n2709, n568, n2017, n5189, n5191, n47,
         n1887, n3539, n2753, n3515, n3794, n3728, n1823, n1210, n4600, n1919,
         n5559, n5958, n5959, n6198, n2573, n1663, n5771, n5766, n6097, n4133,
         n5652, n950, n1132, n4729, n1146, n5150, n954, n5011, n4958, n1021,
         n961, n3922, n2845, n2345, n5501, n966, n1514, n3890, n970, n4842,
         n4841, n973, n974, n4186, n3117, n1902, n3611, n983, n5899, n2055,
         n4938, n2659, n1119, n4006, n6622, n4738, n994, n3640, n1471, n5778,
         n5773, n5827, n5816, n1068, n1651, n3525, n5486, n5485, n5487, n5574,
         n1315, n5680, n1001, n5937, n5936, n6075, n5690, n5692, n5912, n5911,
         n5935, n5502, n5463, n4201, n4200, n2636, n4954, n4955, n4953, n4957,
         n5510, n5480, n5482, n5481, n4378, n4379, n4381, n5908, n5909, n5349,
         n5350, n5224, n5296, n3272, n3271, n3270, n2213, n2212, n2211, n3330,
         n4507, n4617, n4618, n4835, n1251, n3610, n3156, n4688, n4011, n4221,
         n3865, n4132, n4326, n3261, n3830, n5872, n5861, n3719, n3718, n5750,
         n5758, n5752, n3392, n5713, n5703, n5706, n5711, n5709, n5698, n5697,
         n5702, n2420, n1400, n5579, n5580, n1020, n6076, n6074, n6064, n6065,
         n5934, n6112, n6117, n6110, n3615, n1003, n5891, n5890, n5889, n2880,
         n4963, n1161, n1160, n2937, n5537, n5536, n5535, n5538, n5893, n5892,
         n5940, n2833, n4459, n4460, n1005, n6027, n1036, n1007, n4571, n1977,
         n5509, n1681, n1680, n4859, n1250, n5438, n5428, n5175, n6032, n5950,
         n5955, n5517, n5516, n2399, n1255, n1062, n1253, n4663, n2820, n2819,
         n5441, n6037, n4622, n4623, n5340, n2549, n4807, n4141, n2593, n1801,
         n2514, n5527, n2095, n4031, n1057, n4619, n2466, n2569, n2568, n1542,
         n1539, n5422, n3547, n5531, n5530, n5532, n6038, n5953, n5954, n5020,
         n5022, n5080, n4543, n4873, n1884, n4687, n3058, n4530, n4317, n3785,
         n5166, n3803, n3840, n4111, n5387, n6080, n6083, n6009, n6011, n5590,
         n5588, n3725, n5928, n5980, n2864, n5855, n3099, n5732, n5731, n5739,
         n5932, n2863, n5751, n5753, n5755, n1314, n5877, n2976, n5852, n5829,
         n5815, n5806, n5760, n5708, n5705, n5813, n5821, n6084, n6085, n5634,
         n5635, n5576, n5582, n5933, n5575, n5577, n3133, n1307, n6063, n6078,
         n6073, n5971, n5972, n5726, n5696, n5691, n5578, n5581, n5994, n2299,
         n3619, n1289, n1017, n3383, n5215, n2666, n1018, n5704, n4079, n5560,
         n6129, n6130, n6128, n6127, n6126, n6125, n5545, n5543, n5544, n5542,
         n6118, n6116, n1636, n6051, n2881, n2884, n2742, n3410, n6337, n5695,
         n2984, n5664, n5669, n4280, n2286, n6115, n5264, n2497, n6120, n6121,
         n6119, n4202, n6107, n6124, n6113, n6052, n4487, n2805, n1028, n6109,
         n5433, n5431, n5484, n5551, n1032, n6332, n4177, n5352, n3660, n2557,
         n6100, n6099, n6098, n4468, n4462, n4461, n4467, n5943, n5942, n5944,
         n5404, n5941, n5945, n5939, n5511, n5483, n5282, n2663, n3987, n1033,
         n3634, n1034, n5460, n5461, n6103, n6102, n6048, n5029, n4134, n5907,
         n5910, n1335, n1523, n2888, n5285, n5251, n5436, n5435, n3112, n2703,
         n1676, n6041, n6036, n3548, n3766, n4169, n4168, n4170, n5494, n5447,
         n5273, n5271, n5523, n5521, n5956, n5961, n4786, n4041, n1490, n1011,
         n3751, n3017, n3016, n4621, n1040, n4020, n2992, n1252, n3797, n4003,
         n2490, n2528, n4242, n4274, n4516, n4257, n4227, n5269, n5268, n4162,
         n4139, n4140, n5949, n3784, n3783, n6047, n1043, n6046, n3885, n1046,
         n1464, n4451, n1047, n1618, n4126, n6045, n6044, n5283, n1048, n2027,
         n2028, n4032, n1049, n5228, n5225, n1052, n4121, n4123, n6043, n6042,
         n4246, n4237, n4241, n2197, n3888, n2462, n2463, n4936, n1055, n5106,
         n3761, n3971, n1058, n1686, n6096, n6033, n4697, n4698, n3484, n4783,
         n4784, n2885, n5957, n2734, n4846, n1061, n2045, n5409, n2716, n3762,
         n4417, n4321, n5469, n4742, n3795, n5498, n4355, n4922, n4693, n3372,
         n5397, n3849, n4847, n4896, n5904, n4276, n1065, n1256, n2193, n3503,
         n5086, n4886, n1207, n2751, n2029, n3627, n3302, n1089, n1067, n5809,
         n1696, n1072, n1030, n1074, n1073, n2787, n1084, n4616, n2459, n6092,
         n3770, n1664, n1085, n4986, n1086, n1522, n1087, n4881, n1950, n1249,
         n1254, n2571, n3648, n4987, n1235, n1857, n1090, n1092, n3596, n3316,
         n1301, n2022, n2024, n6351, n4739, n2723, n1208, n4002, n1854, n1094,
         n1853, n4685, n2120, n4044, n3322, n1799, n1803, n4500, n2487, n2612,
         n2611, n1097, n3743, n1655, n1485, n3376, n3173, n3174, n3674, n5570,
         n1101, n4433, n5900, n5192, n3773, n4238, n3701, n1106, n2565, n2564,
         n4084, n2595, n4789, n4840, n4156, n4155, n4154, n2896, n2897, n4751,
         n3280, n6326, n1109, n1108, n4951, n2708, n5096, n5095, n5097, n4902,
         n2628, n3909, n5423, n1114, n2058, n1116, n2377, n2376, n1118, n4195,
         n1239, n1121, n3034, n4261, n1125, n1126, n4215, n2186, n2185, n1130,
         n1129, n1128, n4098, n1789, n1131, n1786, n1222, n1303, n1304, n3470,
         n2035, n2036, n4206, n4203, n1135, n5675, n545, n4196, n1770, n4187,
         n1138, n2604, n1139, n1143, n4714, n1144, n6013, n6020, n2592, n3592,
         n711, n2118, n3569, n4374, n2088, n2907, n3297, n4761, n1578, n1165,
         n1580, n1167, n962, n1166, n4696, n4045, n4695, n1168, n2674, n1170,
         n1169, n4858, n1172, n1171, n2392, n1726, n1725, n1174, n6359, n2209,
         n2210, n1173, n1178, n5465, n5503, n5448, n5496, n5495, n3486, n3485,
         n1182, n4918, n1954, n1183, n487, n5033, n3326, n3572, n1186, n2281,
         n1717, n2474, n3714, n3712, n2802, n2026, n4732, n1689, n4728, n1187,
         n1188, n5573, n1608, n5425, n1189, n3488, n3487, n3440, n5426, n3441,
         n1196, n1195, n1192, n4768, n5454, n1198, n2013, n4562, n1199, n2178,
         n1203, n3752, n2979, n2980, n2825, n1205, n1204, n2545, n1209, n1211,
         n4694, n2737, n1213, n1217, n4852, n4844, n4843, n1219, n5948, n4860,
         n1221, n1956, n2349, n2351, n2492, n3411, n1227, n957, n2316, n2978,
         n2312, n1228, n1231, n1229, n2350, n1236, n2001, n6449, n3250, n1555,
         n2244, n1767, n3835, n3837, n3328, n4336, n2413, n2145, n3228, n2678,
         n2679, n4803, n4883, n1242, n2529, n2681, n1244, n1246, n1248, n2192,
         n1795, n6615, n3947, n3626, n3940, n2939, n2898, n2775, n3232, n6193,
         n2713, n3386, n1271, n1045, n5052, n5004, n5005, n1625, n1272, n5003,
         n5054, n1273, n1275, n2177, n969, n1822, n4076, n1377, n6516, n1283,
         n3628, n3106, n3629, n3644, n3643, n3763, n4397, n4398, n2718, n3227,
         n4236, n4482, n4567, n4334, n1547, n1288, n1401, n1291, n1290, n1056,
         n1293, n1292, n3189, n1302, n2080, n1577, n1576, n4709, n2109, n1953,
         n1305, n4879, n4878, n6327, n2171, n2436, n1308, n5681, n1309, n2119,
         n1311, n2665, n2059, n1313, n1312, n5565, n2861, n3819, n3858, n1316,
         n2664, n3518, n2662, n1750, n1317, n1751, n2061, n2060, n3039, n4250,
         n3040, n4672, n1938, n1037, n2661, n4934, n2586, n5028, n2477, n1425,
         n5154, n2655, n5088, n6506, n2037, n1318, n3012, n5160, n1374, n2774,
         n3200, n2931, n3582, n4284, n4299, n3520, n1601, n1923, n3699, n4400,
         n3132, n4877, n46, n4875, n4892, n1325, n1323, n3805, n6203, n1940,
         n3608, n2079, n4910, n2364, n1326, n2822, n1328, n3585, n2008, n2895,
         n2948, n6589, n4828, n1591, n1331, n3066, n1330, n1531, n6459, n1635,
         n2320, n3682, n3681, n3379, n2144, n1334, n2040, n3412, n3345, n2533,
         n3576, n558, n5110, n3151, n1340, n3193, n1341, n3194, n1342, n3198,
         n5362, n3501, n4525, n3195, n3772, n1358, n4218, n1347, n4223, n1349,
         n1348, n2127, n1787, n924, n3143, n3159, n1693, n5794, n3353, n3405,
         n2605, n1353, n1352, n1699, n5257, n3240, n2890, n5258, n1849, n1354,
         n5968, n5927, n5976, n1760, n2419, n1460, n5608, n2986, n5607, n1359,
         n4160, n986, n4083, n3702, n184, n3327, n1364, n1365, n2790, n4508,
         n6617, n1572, n6211, n2372, n2133, n2132, n4273, n5921, n5920, n5925,
         n5781, n1841, n1872, n4458, n440, n4941, n1371, n5622, n4915, n1381,
         n1384, n1386, n2098, n1389, n1388, n2887, n5187, n5186, n1393, n1392,
         n5078, n5146, n5145, n1395, n1399, n1396, n1398, n3111, n5148, n5757,
         n5763, n1402, n1404, n1403, n3889, n3621, n1405, n1409, n5263, n1418,
         n5203, n5152, n2857, n2856, n5202, n1420, n5142, n5204, n5153, n1879,
         n1878, n1426, n1427, n2860, n3374, n2570, n2958, n2441, n1428, n1535,
         n1433, n1513, n1438, n1445, n4808, n1446, n1439, n2030, n1443, n4782,
         n955, n1442, n1441, n1447, n1444, n3352, n1449, n1998, n3335, n4585,
         n1450, n1453, n4004, n1451, n1454, n1456, n4851, n2014, n3546, n1640,
         n6521, n1459, n6210, n3567, n1462, n4799, n4800, n4717, n1466, n1894,
         n2021, n3467, n1508, n1472, n4163, n4164, n2567, n1474, n1473, n1478,
         n1481, n1480, n4937, n4579, n1657, n1656, n1486, n3891, n1487, n3851,
         n1489, n1491, n3748, n1492, n4930, n4929, n1495, n1494, n3897, n1496,
         n2277, n1498, n3899, n1497, n5321, n5767, n2827, n5132, n5129, n5128,
         n5209, n1512, n1743, n1742, n1521, n1519, n1518, n4541, n1526, n4540,
         n1528, n4537, n6605, n4536, n4535, n4893, n3116, n3115, n1532, n5727,
         n3170, n1533, n2579, n2951, n4711, n3222, n3655, n3862, n2100, n4313,
         n1548, n3534, n2432, n2431, n1552, n3993, n1817, n1561, n1558, n1711,
         n3559, n6209, n1560, n4344, n2648, n4629, n1573, n1712, n1574, n2608,
         n1575, n3306, n4403, n1579, n4690, n4948, n2804, n4643, n2150, n2712,
         n1949, n1584, n1588, n1589, n1587, n1590, n2443, n1597, n1604, n2332,
         n1605, n1606, n1614, n1613, n5488, n5434, n1616, n1615, n5464, n3549,
         n1617, n5009, n1624, n4088, n4102, n5214, n5213, n5598, n1631, n6451,
         n2798, n2797, n1642, n3382, n2417, n1643, n2191, n1645, n3243, n3137,
         n1652, n4594, n4591, n1658, n3107, n567, n1659, n1668, n1669, n5534,
         n5533, n1671, n1670, n4773, n4772, n5915, n5917, n5914, n1677, n1679,
         n5411, n1682, n4268, n4269, n1688, n3428, n3321, n2903, n3168, n2266,
         n1695, n1697, n2955, n2891, n5207, n5261, n5262, n5309, n4700, n1703,
         n4702, n1704, n1706, n1705, n1708, n1707, n4419, n4420, n4421, n3314,
         n2624, n4978, n6520, n2942, n1718, n2947, n2998, n1722, n5353, n2062,
         n2656, n4787, n1732, n1731, n1730, n1734, n1738, n1737, n1736, n1740,
         n1888, n3402, n6330, n4477, n2365, n1757, n1758, n1763, n5473, n1761,
         n1762, n1766, n6619, n2279, n4116, n4114, n1771, n4109, n2273, n4208,
         n4082, n2335, n2352, n3449, n4757, n4756, n4755, n4710, n1793, n1792,
         n2190, n2590, n1797, n1796, n5062, n1802, n5018, n5016, n1816, n1815,
         n1809, n1806, n6303, n1814, n1811, n1818, n1821, n1819, n2033, n2990,
         n3229, n4052, n4053, n4054, n1838, n4464, n1843, n4068, n2765, n6329,
         n1951, n1856, n1855, n1859, n1861, n1860, n987, n3169, n1866, n6602,
         n2034, n5001, n5000, n5122, n5123, n2356, n3574, n3093, n3429, n3510,
         n3358, n1883, n3312, n6263, n1936, n1889, n1890, n4036, n4035, n1891,
         n3956, n4043, n1892, n2002, n1895, n4560, n1896, n6104, n4255, n1899,
         n4253, n3612, n5974, n5979, n1904, n1906, n2677, n3341, n6381, n5662,
         n5663, n1916, n1922, n3812, n3997, n3711, n1926, n1924, n1931, n3577,
         n4940, n5109, n6460, n5064, n1939, n4572, n2680, n1959, n1958, n4744,
         n5130, n3109, n1967, n1966, n1965, n1970, n1968, n3965, n6251, n3925,
         n2996, n5048, n2764, n3630, n2115, n189, n3216, n3079, n2577, n4415,
         n5219, n1989, n2727, n2472, n4745, n4836, n4949, n4950, n3908, n3906,
         n6588, n2000, n6357, n5859, n5325, n5327, n4644, n4639, n2007, n2531,
         n3152, n4503, n3439, n4638, n2016, n2015, n4081, n3729, n4492, n4493,
         n4588, n4659, n4129, n2582, n2446, n2020, n2632, n2631, n2801, n2800,
         n4191, n4190, n2041, n3255, n5012, n3669, n3532, n2047, n3531, n2046,
         n5081, n5082, n2814, n2053, n3599, n2052, n2817, n2057, n2739, n5371,
         n5290, n3558, n5492, n2067, n5567, n2068, n2071, n2070, n3028, n3027,
         n2075, n5114, n5116, n4996, n5083, n2078, n5195, n3230, n4491, n6344,
         n3347, n2105, n2106, n2317, n2761, n2763, n2112, n4278, n2428, n2429,
         n2675, n2123, n2121, n3739, n3740, n3671, n2139, n2138, n6155, n2142,
         n2149, n4325, n2158, n2402, n2160, n4324, n2162, n2667, n2165, n4646,
         n2164, n2169, n2714, n3223, n3841, n2706, n3649, n3796, n3798, n3786,
         n4249, n3035, n965, n2427, n6293, n2271, n4213, n2194, n2203, n2204,
         n2207, n2206, n3697, n5247, n3423, n958, n3301, n3857, n2214, n3859,
         n3821, n3822, n2217, n2216, n3293, n4359, n6455, n4444, n4033, n6191,
         n2224, n2225, n2228, n2227, n2232, n4148, n5657, n2233, n2234, n5648,
         n5649, n5650, n3274, n2236, n2293, n3732, n2237, n5733, n4305, n3212,
         n2240, n3356, n2450, n2449, n4181, n4180, n2250, n2252, n2260, n2259,
         n2258, n3183, n3186, n3910, n2263, n4119, n4120, n2264, n5746, n2265,
         n5741, n5728, n5783, n5784, n5797, n5796, n5802, n2269, n5599, n2705,
         n3471, n3498, n5380, n5379, n5625, n5382, n3380, n2282, n2777, n3381,
         n2284, n3848, n2288, n2287, n2862, n6133, n6131, n5938, n2338, n5372,
         n4157, n2341, n2340, n5550, n2344, n2342, n5497, n2343, n5346, n5348,
         n5549, n3508, n2346, n3451, n2359, n2361, n2362, n3690, n2363, n6180,
         n5710, n5715, n3041, n4820, n4819, n2370, n3556, n2379, n2378, n4544,
         n5182, n2953, n5178, n3673, n2380, n5181, n2381, n5098, n3295, n3119,
         n991, n2387, n2385, n4008, n2390, n3398, n2575, n2395, n2394, n5063,
         n5066, n2396, n5319, n2400, n3413, n3334, n5226, n5229, n2404, n2407,
         n3688, n3686, n2414, n5037, n2425, n4270, n2433, n2455, n2454, n2456,
         n4620, n2475, n2476, n2482, n2493, n3360, n5977, n5318, n2494, n2495,
         n2499, n5265, n2496, n2501, n2504, n2982, n2505, n6012, n2981, n5057,
         n5440, n5061, n5561, n2521, n5370, n6508, n5367, n2525, n2527, n5823,
         n3978, n3977, n5410, n6524, n4898, n5396, n5467, n5179, n3357, n2553,
         n2554, n5280, n2558, n5356, n3661, n2555, n2556, n5351, n2560, n5281,
         n5279, n6239, n2673, n5316, n5597, n3397, n5337, n4634, n3104, n2584,
         n2585, n3092, n3091, n2598, n2606, n2610, n2609, n2616, n2615, n2618,
         n2617, n2620, n2619, n2911, n2621, n2625, n2626, n2627, n3252, n4884,
         n2634, n4345, n2650, n5087, n5284, n2660, n3517, n3963, n3633, n2670,
         n2671, n2672, n3689, n565, n2686, n2684, n2685, n2687, n4010, n2697,
         n2696, n2698, n4494, n3187, n3597, n5104, n3505, n953, n5221, n5222,
         n3320, n4252, n6040, n6034, n2988, n4310, n5814, n5824, n6453, n3098,
         n4678, n4673, n4676, n3472, n6457, n3652, n3128, n4832, n3445, n2915,
         n3490, n5445, n3781, n3566, n4448, n4440, n5121, n5067, n5068, n3309,
         n4204, n6178, n4383, n4386, n5499, n4101, n4096, n4645, n5960, n6123,
         n6105, n4260, n4263, n6201, n4264, n6376, n2938, n3005, n2782, n2780,
         n5981, n6066, n6067, n6108, n4125, n4127, n5651, n5654, n5656, n5659,
         n5655, n4117, n4112, n5693, n4234, n4233, n5712, n5714, n5775, n5747,
         n5744, n6522, n5748, n5743, n5754, n5799, n5800, n5791, n5803, n5837,
         n5849, n5605, n5606, n6025, n5963, n2851, n5966, n5964, n4813, n3639,
         n3878, n2730, n3071, n3437, n4675, n3246, n4944, n3653, n3969, n3343,
         n3054, n3053, n4062, n4429, n4825, n4827, n3442, n5398, n3543, n4590,
         n3964, n2866, n2867, n4453, n2919, n4454, n3177, n4021, n5249, n5278,
         n5442, n4897, n5466, n5363, n5415, n5407, n5339, n3443, n5208, n5211,
         n5347, n5896, n426, n3847, n3846, n3007, n4980, n5522, n5520, n6077,
         n4110, n5688, n3416, n6505, n3414, n5858, n5600, n6661, n5333, n6509,
         n2711, n6114, n5831, n3387, n3721, n3717, n3716, n5850, n3715, n6006,
         n5998, n6008, n6004, n6007, n6003, n6072, n6002, n5878, n5879, n5583,
         n5586, n6137, n5646, n5645, n5644, n5653, n5661, n5668, n5666, n5674,
         n5673, n5679, n5701, n5700, n5801, n5811, n5812, n5810, n2702, n2704,
         n2710, n4522, n5432, n5540, n2725, n2726, n2729, n2732, n2740, n2745,
         n2747, n5025, n3399, n3311, n2754, n2759, n2760, n5046, n2762, n5050,
         n5394, n2768, n4956, n2772, n4533, n2781, n2778, n3390, n5842, n5624,
         n5375, n5623, n4971, n2793, n2794, n2795, n4947, n2807, n5601, n5993,
         n5992, n4060, n2815, n2816, n3142, n5476, n2829, n3288, n2832, n3391,
         n5887, n289, n4719, n3605, n2841, n4603, n2842, n4602, n2844, n2850,
         n6111, n2908, n5141, n5140, n2858, n2859, n5135, n2875, n2873, n6071,
         n5612, n6526, n4988, n2886, n4647, n5628, n5969, n5603, n5604, n5233,
         n5234, n6328, n4815, n6095, n2892, n2893, n2894, n6094, n5161, n5162,
         n5163, n5723, n5724, n2294, n5719, n6199, n2900, n6001, n5584, n5591,
         n5871, n5602, n5631, n5378, n6447, n3001, n2906, n3310, n3432, n6185,
         n6616, n3992, n5420, n3424, n3464, n4793, n4013, n3004, n4521, n4574,
         n2935, n2934, n5385, n2941, n2940, n4553, n2944, n2943, n2946, n3287,
         n2959, n3541, n5793, n2970, n3914, n4428, n4427, n2985, n4984, n4983,
         n997, n4985, n2991, n4018, n4016, n4017, n2994, n3495, n3000, n2999,
         n3203, n3006, n3014, n4625, n6570, n3018, n4384, n3019, n6528, n4337,
         n4026, n3031, n3030, n4259, n4265, n3036, n3037, n3038, n3349, n579,
         n3043, n3045, n3044, n3960, n3047, n3046, n3962, n3048, n3055, n4471,
         n4343, n3081, n3084, n3578, n3579, n3097, n3102, n3101, n3406, n5856,
         n3100, n5857, n3560, n3120, n5860, n3377, n3378, n3317, n3135, n3138,
         n3139, n3141, n3140, n3144, n3145, n4885, n4595, n4596, n6213, n3146,
         n3148, n3363, n5682, n6138, n6136, n3790, n3163, n3162, n3164, n3678,
         n5627, n3676, n3167, n3276, n3180, n3179, n3181, n4597, n3182, n1100,
         n5507, n4226, n5193, n5194, n5137, n5138, n945, n3226, n4039, n3233,
         n5843, n5848, n2736, n4870, n3254, n4857, n3269, n5030, n3749, n3279,
         n3277, n4627, n4292, n4925, n5841, n3340, n3339, n6156, n5528, n3354,
         n5847, n5846, n3361, n5685, n3366, n4358, n3373, n3601, n4887, n3394,
         n4357, n908, n3401, n3400, n3789, n3422, n3419, n3425, n4943, n5015,
         n3614, n3433, n3444, n5468, n3455, n185, n3454, n4182, n4230, n3459,
         n3460, n4312, n3497, n3921, n4891, n5462, n3489, n3737, n3499, n3506,
         n4377, n3513, n3514, n5232, n3519, n5830, n4707, n3544, n3542, n5417,
         n1015, n5845, n4235, n3998, n3565, n4029, n4028, n3618, n4283, n3590,
         n4089, n4166, n4225, n4165, n3799, n2733, n3632, n3637, n3638, n3884,
         n3651, n344, n5922, n6350, n5313, n5026, n3677, n3679, n4209, n4207,
         n5990, n5595, n5594, n3687, n3771, n5180, n5250, n3698, n3720, n6360,
         n5874, n5310, n6018, n4587, n4328, n4329, n3735, n3734, n3741, n3750,
         n3754, n6464, n5785, n5786, n5787, n5832, n4981, n2878, n5965, n4665,
         n3765, n5587, n5585, n3768, n4725, n4679, n4790, n4831, n5267, n4446,
         n4449, n4439, n3788, n5124, n5272, n5270, n2756, n5157, n4128, n5854,
         n5978, n5779, n3780, n3782, n4092, n4823, n3787, n3791, n3793, n3808,
         n3810, n3818, n5101, n3829, n3839, n3850, n4609, n3874, n3873, n3875,
         n3876, n3879, n3893, n3929, n3918, n762, n3951, n3970, n3972, n3973,
         n3989, n3995, n4014, n4022, n4023, n4024, n4030, n4047, n4049, n4063,
         n4066, n4093, n4094, n4113, n4122, n4136, n4147, n4146, n4153, n4178,
         n4210, n4220, n4222, n4258, n4256, n4240, n4251, n4262, n4286, n4290,
         n4311, n6026, n4361, n4364, n4362, n4367, n4380, n4391, n4390, n4396,
         n4393, n4395, n4399, n4027, n4425, n4426, n4424, n4423, n4431, n4438,
         n4441, n4495, n4532, n4547, n4548, n4561, n4613, n4610, n4615, n4660,
         n4664, n4680, n4682, n4699, n4706, n4722, n6406, n4727, n4792, n4806,
         n4809, n6182, n4818, n4817, n4822, n4830, n4848, n4850, n4849, n6458,
         n4926, n4932, n946, n4945, n4990, n4992, n4991, n4993, n5007, n5006,
         n6153, n5071, n610, n5100, n5103, n5102, n5107, n5165, n5125, n5159,
         n5158, n5199, n5196, n5198, n5223, n6674, n5230, n5227, n5236, n5237,
         n5245, n5243, n5244, n888, n5256, n6424, n5254, n5274, n6154, n5338,
         n5344, n5343, n5366, n5399, n5403, n5401, n5400, n5402, n5408, n5406,
         n5405, n5416, n5539, n5430, n5419, n5429, n5421, n5443, n5444, n5446,
         n5456, n5500, n5470, n5475, n5474, n5479, n5478, n5512, n5548, n5515,
         n5519, n5518, n5524, n5906, n5569, n5589, n5885, n5614, n5615, n5613,
         n5619, n5638, n5637, n6056, n5636, n5639, n5641, n5640, n5683, n325,
         n5684, n5687, n5720, n5737, n5736, n5738, n5740, n5756, n5749, n5759,
         n5762, n5761, n5770, n5805, n3427, n6375, n5820, n5826, n5833, n5882,
         n5880, n5881, n5898, n5903, n5902, n6585, n5901, n5905, n5946, n5962,
         n6058, n5967, n5985, n5988, n6101, n6057, n6060, n6061, n6069, n6166,
         n3767, n6082, n496, n6091, n6087, n6088, n6089, n6090, n6106, n295,
         n209, n6165, n28, n4456, n4455, n6413, n4970, n3256, n848, n1568,
         n1567, n4445, n138, n151, n3210, n4766, n3512, n85, n1463, n3968,
         n4330, n2965, n5923, n1367, n4086, n396, n2484, n2485, n4418, n4497,
         n872, n352, n3685, n3665, n469, n193, n814, n2997, n6495, n2701,
         n5643, n5002, n5642, n3022, n704, n4791, n379, n19, n3623, n4352,
         n3804, n4385, n956, n1537, n1536, n316, n3057, n5017, n355, n4243,
         n3967, n4198, n2011, n3926, n273, n447, n1122, n905, n1900, n1901,
         n6054, n768, n3946, n5686, n834, n5730, n6423, n6348, n5825, n6194,
         n5632, n1232, n5365, n5231, n2247, n4771, n3616, n1488, n1053, n776,
         n497, n3281, n632, n1804, n1499, n6378, n64, n4546, n3507, n2792,
         n2175, n2174, n1975, n3668, n6342, n6343, n4306, n5790, n6164, n806,
         n6171, n2292, n2901, n6405, n2122, n2574, n5126, n6339, n6338, n6253,
         n4712, n6229, n1592, n2552, n1416, n1415, n3707, n3231, n6333, n128,
         n1269, n6371, n6372, n6374, n634, n631, n1632, n6361, n6368, n6316,
         n6448, n6237, n4341, n1839, n6390, n3493, n4366, n6181, n6159, n4797,
         n6184, n3300, n1784, n3299, n350, n6172, n6170, n2439, n5455, n859,
         n6162, n1026, n6163, n1764, n6363, n6297, n3332, n6169, n2838, n2012,
         n6173, n6345, n6174, n1527, n1414, n1837, n4301, n2285, n6175, n6176,
         n6177, n4171, n6618, n6179, n4224, n6264, n3666, n6188, n2905, n6189,
         n4716, n4422, n1069, n2977, n1298, n1264, n3826, n1690, n2422, n6212,
         n6216, n6220, n6219, n6222, n6223, n2416, n1807, n2418, n6224, n6226,
         n6225, n6291, n6228, n226, n225, n3319, n6256, n6422, n3477, n6230,
         n4931, n6231, n6232, n269, n4294, n6233, n6235, n6234, n3948, n6236,
         n6157, n4173, n2056, n6238, n6240, n6241, n6245, n6243, n6242, n6246,
         n6249, n429, n1541, n6250, n6252, n6437, n6436, n6254, n6403, n5085,
         n6255, n6385, n6258, n4804, n6260, n6259, n4303, n3384, n5259, n6265,
         n6439, n6266, n439, n3033, n2614, n6267, n4518, n5156, n4108, n428,
         n1366, n6268, n122, n6269, n495, n6270, n6272, n6274, n6273, n6276,
         n6275, n2452, n6277, n97, n2635, n3026, n6590, n6468, n6278, n3094,
         n6279, n6283, n5864, n6284, n2623, n2622, n6286, n6287, n191, n692,
         n6289, n6290, n3777, n6294, n6295, n1184, n6296, n2572, n6298, n6365,
         n451, n6299, n1357, n6601, n1915, n876, n1111, n335, n2447, n6300,
         n287, n6302, n6301, n1525, n1921, n4103, n6304, n6418, n6305, n6306,
         n6404, n6307, n6407, n6308, n6309, n3902, n3021, n2126, n6310, n3436,
         n6431, n6311, n2993, n364, n6315, n4368, n3067, n6317, n5115, n6319,
         n6318, n6320, n5304, n6321, n6322, n2904, n3709, n6474, n3298, n3134,
         n835, n590, n3604, n4371, n4199, n6334, n774, n3294, n5164, n3845,
         n886, n6340, n6341, n6346, n6347, n4928, n2776, n4436, n1948, n6349,
         n2532, n5093, n6352, n6353, n6355, n6354, n6356, n2478, n3920, n1286,
         n942, n6358, n3844, n6362, n6364, n6369, n6367, n6370, n6373, n6379,
         n6432, n6380, n6382, n6384, n6383, n2652, n6386, n6388, n6387, n1990,
         n6392, n6393, n3550, n1278, n1563, n6394, n6395, n6397, n6398, n6399,
         n2136, n2134, n6401, n6400, n4360, n3103, n2924, n2535, n1078, n1987,
         n456, n6408, n1115, n6410, n6411, n187, n6412, n6415, n6530, n6417,
         n6419, n6420, n6421, n1952, n6425, n6427, n6426, n6465, n6428, n6433,
         n6434, n6435, n1156, n2091, n2591, n6438, n6442, n6443, n3667, n6444,
         n3260, n639, n1262, n4432, n6621, n207, n5205, n1103, n2318, n2536,
         n1666, n6288, n1070, n904, n3483, n623, n399, n680, n6492, n4658,
         n4167, n2855, n6227, n291, n2509, n570, n1662, n302, n5505, n2854,
         n6192, n2481, n4683, n901, n879, n3171, n250, n1897, n5735, n5844,
         n2771, n3123, n1566, n797, n577, n2220, n798, n4347, n3225, n1945,
         n310, n35, n312, n313, n4501, n2486, n1220, n2503, n6414, n2464,
         n6167, n6053, n6049, n1654, n6257, n6604, n4648, n6491, n6613, n2728,
         n2147, n2507, n4104, n5504, n6606, n3759, n152, n6593, n1691, n1692,
         n1452, n6658, n6132, n5108, n5626, n3375, n6461, n2551, n6440, n6649,
         n6469, n6597, n6507, n6285, n3692, n6566, n6479, n938, n6620, n6488,
         n1382, n6680, n6462, n6463, n6466, n6467, n3641, n2141, n6578, n6470,
         n5395, n5328, n6471, n6482, n6472, n6473, n6581, n6475, n2222, n6477,
         n6476, n6168, n6496, n6478, n6480, n963, n6656, n533, n578, n6481,
         n2221, n6561, n3122, n1893, n6483, n5618, n6626, n6625, n6484, n6281,
         n6486, n6485, n6533, n4927, n1319, n6487, n131, n6489, n3185, n3744,
         n6640, n6490, n5863, n6010, n6639, n6493, n6494, n5329, n6672, n6628,
         n3662, n4074, n6497, n6498, n2722, n2542, n6499, n6500, n6592, n6501,
         n6503, n6502, n6552, n2960, n6510, n4960, n6512, n6550, n6517, n6518,
         n6523, n3199, n6531, n6536, n6532, n6644, n4718, n6534, n6535, n6537,
         n6538, n6539, n6540, n6541, n6635, n6542, n6591, n6543, n6545, n6544,
         n6547, n6546, n6572, n6669, n6548, n3564, n6549, n6551, n899, n6553,
         n6555, n6554, n6556, n6557, n6559, n6560, n6563, n6562, n6564, n57,
         n6565, n6568, n6567, n6668, n6571, n6574, n6573, n6576, n6575, n3511,
         n6577, n6664, n6663, n6579, n996, n6580, n6611, n6582, n6583, n6584,
         n6650, n6586, n2018, n6594, n6595, n2257, n6599, n6598, n6600, n6603,
         n906, n2125, n6612, n6645, n3880, n4291, n6629, n6627, n6630, n6633,
         n6634, n6638, n5865, n5866, n669, n5312, n6636, n6637, n6641, n6642,
         n6643, n6647, n6646, n6135, n6648, n6651, n6652, n6653, n6657, n6660,
         n6659, n2301, n6662, n968, n6665, n6666, n6667, n6675, n6671, n6670,
         n6673, n6676, n6677, n6678, n6679, n1476, n1475, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6694,
         n6695, n6696, n4750, n6697, n6698, n3583, n6699;

  BUF_X4 U2 ( .A(n5798), .Z(n976) );
  NAND2_X2 U3 ( .A1(n5808), .A2(n5807), .ZN(n5838) );
  NOR2_X2 U4 ( .A1(n2157), .A2(n5918), .ZN(n4973) );
  NAND2_X2 U5 ( .A1(n5610), .A2(n5609), .ZN(n369) );
  NAND2_X2 U7 ( .A1(n1243), .A2(n989), .ZN(n4583) );
  NAND2_X2 U10 ( .A1(n1634), .A2(n5036), .ZN(n5091) );
  NAND2_X2 U12 ( .A1(n1756), .A2(n1755), .ZN(n3125) );
  INV_X4 U13 ( .A(n690), .ZN(n3409) );
  NAND2_X2 U15 ( .A1(n520), .A2(n521), .ZN(n4907) );
  NOR2_X2 U18 ( .A1(n4281), .A2(n4282), .ZN(n2114) );
  NAND2_X2 U19 ( .A1(n3158), .A2(n5357), .ZN(n5556) );
  NAND2_X2 U21 ( .A1(n1150), .A2(n1152), .ZN(n5694) );
  NAND2_X2 U23 ( .A1(n3245), .A2(n3248), .ZN(n4906) );
  NAND2_X2 U25 ( .A1(n604), .A2(n605), .ZN(n3561) );
  NOR2_X2 U26 ( .A1(n3421), .A2(n3824), .ZN(n3823) );
  NAND2_X2 U27 ( .A1(n2170), .A2(n2523), .ZN(n3023) );
  NAND2_X2 U28 ( .A1(n1863), .A2(n1862), .ZN(n2201) );
  NAND2_X2 U30 ( .A1(n811), .A2(n812), .ZN(n557) );
  NAND2_X2 U34 ( .A1(n5359), .A2(n5358), .ZN(n5457) );
  NAND2_X2 U35 ( .A1(n3237), .A2(n3475), .ZN(n3747) );
  NOR2_X2 U38 ( .A1(n5079), .A2(n3540), .ZN(n1225) );
  NOR2_X2 U39 ( .A1(n2871), .A2(n2874), .ZN(n2870) );
  NAND2_X2 U40 ( .A1(n3251), .A2(n4741), .ZN(n2314) );
  NAND2_X2 U41 ( .A1(n2103), .A2(n4743), .ZN(n1960) );
  NAND2_X2 U44 ( .A1(n1193), .A2(n3217), .ZN(n1397) );
  NAND2_X2 U46 ( .A1(n1646), .A2(n1647), .ZN(n2076) );
  NOR3_X2 U50 ( .A1(n463), .A2(n464), .A3(n2836), .ZN(n461) );
  NOR2_X1 U51 ( .A1(n2828), .A2(n3915), .ZN(n3916) );
  INV_X2 U52 ( .A(n159), .ZN(n1477) );
  NOR2_X2 U54 ( .A1(n3404), .A2(n4692), .ZN(n4762) );
  NOR2_X2 U58 ( .A1(n5075), .A2(n947), .ZN(n1646) );
  NAND2_X2 U61 ( .A1(n3242), .A2(n3241), .ZN(n5167) );
  INV_X4 U63 ( .A(n4239), .ZN(n4217) );
  NOR2_X2 U68 ( .A1(n5079), .A2(n4788), .ZN(n2596) );
  NAND2_X2 U70 ( .A1(b[0]), .A2(n1287), .ZN(n4100) );
  NOR3_X2 U71 ( .A1(n923), .A2(n3435), .A3(n1554), .ZN(n921) );
  NAND2_X2 U73 ( .A1(a[23]), .A2(b[12]), .ZN(n5294) );
  NOR2_X1 U74 ( .A1(n5190), .A2(n3760), .ZN(n4607) );
  INV_X2 U75 ( .A(b[11]), .ZN(n865) );
  INV_X4 U78 ( .A(n3533), .ZN(n3642) );
  NOR2_X2 U80 ( .A1(n4770), .A2(n3617), .ZN(n3324) );
  NAND2_X2 U81 ( .A1(n2717), .A2(n3562), .ZN(n2270) );
  NAND2_X2 U82 ( .A1(n1147), .A2(b[10]), .ZN(n4489) );
  NAND2_X2 U88 ( .A1(n3757), .A2(a[0]), .ZN(n3209) );
  INV_X4 U93 ( .A(n5477), .ZN(n5947) );
  INV_X4 U96 ( .A(b[15]), .ZN(n984) );
  INV_X4 U98 ( .A(n4677), .ZN(n1064) );
  INV_X4 U99 ( .A(n29), .ZN(n1194) );
  NOR2_X2 U103 ( .A1(a[1]), .A2(a[2]), .ZN(n635) );
  INV_X4 U106 ( .A(b[11]), .ZN(n981) );
  NOR2_X2 U108 ( .A1(n513), .A2(b[19]), .ZN(n1329) );
  NAND2_X2 U112 ( .A1(a[3]), .A2(a[4]), .ZN(n734) );
  NAND2_X4 U124 ( .A1(a[13]), .A2(a[14]), .ZN(n3952) );
  NAND2_X2 U126 ( .A1(n4733), .A2(n753), .ZN(n3220) );
  NAND2_X2 U127 ( .A1(n1847), .A2(n5293), .ZN(n2412) );
  NAND2_X4 U128 ( .A1(n194), .A2(n911), .ZN(n5718) );
  NAND2_X2 U129 ( .A1(n2305), .A2(n304), .ZN(n614) );
  NOR2_X4 U130 ( .A1(n5413), .A2(n5412), .ZN(n5541) );
  INV_X4 U131 ( .A(n5541), .ZN(n5414) );
  NAND2_X2 U137 ( .A1(n2043), .A2(n4952), .ZN(n808) );
  XNOR2_X2 U138 ( .A(n2093), .B(n949), .ZN(n1633) );
  NAND2_X2 U139 ( .A1(n5514), .A2(n5513), .ZN(n5547) );
  NOR2_X2 U141 ( .A1(n5235), .A2(b[23]), .ZN(n2914) );
  XOR2_X2 U142 ( .A(a[3]), .B(b[16]), .Z(n2744) );
  XOR2_X2 U146 ( .A(a[3]), .B(b[14]), .Z(n2715) );
  NOR2_X4 U147 ( .A1(a[3]), .A2(a[1]), .ZN(n4834) );
  NAND2_X1 U151 ( .A1(n5074), .A2(n5951), .ZN(n2116) );
  NOR2_X2 U152 ( .A1(n5074), .A2(b[5]), .ZN(n2309) );
  OAI21_X1 U155 ( .B1(n2786), .B2(n2933), .A(n5376), .ZN(n2785) );
  INV_X4 U159 ( .A(n5119), .ZN(n5117) );
  OAI21_X1 U160 ( .B1(n5197), .B2(a[15]), .A(b[8]), .ZN(n1981) );
  INV_X8 U161 ( .A(a[13]), .ZN(n3369) );
  NAND2_X4 U164 ( .A1(n529), .A2(n528), .ZN(n6093) );
  NOR2_X2 U168 ( .A1(n2700), .A2(n4777), .ZN(n2256) );
  OAI21_X2 U169 ( .B1(n3882), .B2(n2700), .A(n3881), .ZN(n3883) );
  NAND2_X2 U171 ( .A1(n328), .A2(n4559), .ZN(n1) );
  NAND2_X2 U173 ( .A1(n2), .A2(n394), .ZN(n1411) );
  NAND2_X2 U174 ( .A1(n392), .A2(n5300), .ZN(n2) );
  XNOR2_X2 U175 ( .A(n3), .B(n3823), .ZN(n3985) );
  XNOR2_X2 U176 ( .A(n3813), .B(n3814), .ZN(n3) );
  NAND2_X2 U178 ( .A1(n4), .A2(n391), .ZN(n1406) );
  NAND2_X2 U180 ( .A1(n5184), .A2(n564), .ZN(n5185) );
  AOI21_X2 U181 ( .B1(n5242), .B2(n5241), .A(n5240), .ZN(n5303) );
  NOR2_X2 U182 ( .A1(n5169), .A2(n5), .ZN(n5242) );
  INV_X2 U183 ( .A(n6), .ZN(n5) );
  NAND2_X2 U184 ( .A1(n5168), .A2(n1999), .ZN(n6) );
  NAND2_X2 U185 ( .A1(n1429), .A2(n1430), .ZN(n283) );
  NAND2_X2 U186 ( .A1(n1534), .A2(n2189), .ZN(n1429) );
  NOR2_X2 U187 ( .A1(n4733), .A2(n753), .ZN(n3149) );
  INV_X2 U189 ( .A(n4480), .ZN(n7) );
  NAND2_X2 U191 ( .A1(n8), .A2(n1093), .ZN(n170) );
  NAND2_X2 U192 ( .A1(n2184), .A2(n4463), .ZN(n8) );
  NAND2_X4 U195 ( .A1(n1852), .A2(n2548), .ZN(n3755) );
  INV_X4 U196 ( .A(n3755), .ZN(n1851) );
  NAND2_X2 U197 ( .A1(n1408), .A2(n971), .ZN(n1407) );
  INV_X4 U203 ( .A(n5308), .ZN(n1019) );
  NAND3_X2 U205 ( .A1(n2430), .A2(n2274), .A3(n2275), .ZN(n2137) );
  NOR2_X2 U206 ( .A1(n1193), .A2(b[2]), .ZN(n4051) );
  OAI22_X2 U209 ( .A1(n4118), .A2(n4490), .B1(b[3]), .B2(n6183), .ZN(n4142) );
  NAND2_X2 U214 ( .A1(n3856), .A2(n3855), .ZN(n3898) );
  NAND3_X2 U215 ( .A1(n3730), .A2(n4333), .A3(n4332), .ZN(n2124) );
  XNOR2_X2 U217 ( .A(n11), .B(n4450), .ZN(n3042) );
  NAND2_X2 U222 ( .A1(n14), .A2(n13), .ZN(n1756) );
  NAND2_X2 U224 ( .A1(n6149), .A2(n4472), .ZN(n14) );
  NAND2_X2 U225 ( .A1(n3265), .A2(n909), .ZN(n4527) );
  NOR2_X2 U228 ( .A1(n251), .A2(n3957), .ZN(n4034) );
  NAND2_X2 U229 ( .A1(n3894), .A2(n1050), .ZN(n1432) );
  NAND2_X2 U230 ( .A1(n261), .A2(n262), .ZN(n264) );
  NOR2_X2 U232 ( .A1(n3049), .A2(n3050), .ZN(n15) );
  NAND2_X2 U233 ( .A1(n3369), .A2(b[7]), .ZN(n4363) );
  BUF_X4 U235 ( .A(n2009), .Z(n16) );
  NAND2_X2 U237 ( .A1(n174), .A2(n941), .ZN(n1583) );
  NAND2_X4 U240 ( .A1(n2909), .A2(n2910), .ZN(n2912) );
  AOI21_X2 U241 ( .B1(n6336), .B2(n5834), .A(n2006), .ZN(n5323) );
  AOI22_X2 U244 ( .A1(n1051), .A2(n1225), .B1(n2104), .B2(n3802), .ZN(n17) );
  NAND2_X2 U246 ( .A1(n3694), .A2(n3693), .ZN(n3307) );
  NOR2_X2 U248 ( .A1(n2187), .A2(n1363), .ZN(n1362) );
  NAND2_X2 U250 ( .A1(n1973), .A2(n4496), .ZN(n2511) );
  NAND2_X2 U251 ( .A1(n2868), .A2(n2869), .ZN(n4496) );
  INV_X4 U255 ( .A(n4478), .ZN(n3446) );
  INV_X4 U256 ( .A(n2566), .ZN(n4085) );
  NAND2_X2 U257 ( .A1(n813), .A2(n16), .ZN(n816) );
  AOI22_X2 U258 ( .A1(n4350), .A2(n4351), .B1(n4349), .B2(n3308), .ZN(n4354)
         );
  NAND2_X2 U259 ( .A1(n21), .A2(n20), .ZN(n3072) );
  NAND2_X2 U261 ( .A1(n4405), .A2(b[17]), .ZN(n21) );
  INV_X4 U267 ( .A(n2411), .ZN(n674) );
  NAND2_X2 U268 ( .A1(n22), .A2(n323), .ZN(n3234) );
  NAND2_X2 U269 ( .A1(n321), .A2(n4566), .ZN(n22) );
  NAND2_X2 U272 ( .A1(n4267), .A2(n4266), .ZN(n5699) );
  NAND2_X2 U274 ( .A1(n23), .A2(n288), .ZN(n4254) );
  NAND2_X2 U276 ( .A1(n1582), .A2(n1581), .ZN(n4557) );
  INV_X2 U280 ( .A(n24), .ZN(\d[15]_BAR ) );
  NOR2_X2 U281 ( .A1(n27), .A2(n25), .ZN(n24) );
  NOR2_X2 U284 ( .A1(n5776), .A2(n5774), .ZN(n27) );
  NOR2_X2 U285 ( .A1(n6454), .A2(n771), .ZN(n5725) );
  NAND2_X2 U287 ( .A1(n2031), .A2(n4565), .ZN(n323) );
  INV_X2 U296 ( .A(n760), .ZN(n29) );
  BUF_X4 U297 ( .A(n4734), .Z(n30) );
  NAND2_X1 U298 ( .A1(n1571), .A2(n3283), .ZN(n651) );
  XNOR2_X2 U299 ( .A(n2283), .B(n4734), .ZN(n1571) );
  INV_X4 U300 ( .A(n3468), .ZN(n1470) );
  NAND2_X2 U301 ( .A1(n4319), .A2(n4318), .ZN(n2676) );
  NAND3_X2 U302 ( .A1(n1008), .A2(n1152), .A3(n6187), .ZN(n1117) );
  NAND2_X4 U304 ( .A1(n2229), .A2(n31), .ZN(n4636) );
  NAND3_X2 U305 ( .A1(n3446), .A2(n2375), .A3(n6366), .ZN(n31) );
  NAND2_X2 U308 ( .A1(n3069), .A2(n3070), .ZN(n4040) );
  NAND2_X2 U310 ( .A1(n3197), .A2(n3196), .ZN(n1831) );
  NAND2_X2 U312 ( .A1(n869), .A2(n868), .ZN(n5629) );
  NAND2_X2 U313 ( .A1(n2003), .A2(n584), .ZN(n1469) );
  NAND2_X2 U315 ( .A1(n3753), .A2(n3645), .ZN(n2215) );
  INV_X2 U318 ( .A(n1700), .ZN(n866) );
  NAND2_X2 U319 ( .A1(n1702), .A2(n1701), .ZN(n1700) );
  INV_X4 U320 ( .A(n4465), .ZN(n1093) );
  NAND2_X2 U323 ( .A1(n32), .A2(n444), .ZN(n1333) );
  NAND2_X2 U324 ( .A1(n442), .A2(n443), .ZN(n32) );
  NAND2_X2 U325 ( .A1(n1483), .A2(n1482), .ZN(n633) );
  NAND2_X2 U326 ( .A1(n5252), .A2(n2291), .ZN(n871) );
  NAND2_X2 U327 ( .A1(n4061), .A2(n4055), .ZN(n4057) );
  NAND2_X4 U328 ( .A1(n4601), .A2(b[20]), .ZN(n3606) );
  AOI21_X2 U329 ( .B1(n5188), .B2(n1394), .A(n1390), .ZN(n5239) );
  NOR2_X4 U330 ( .A1(n1391), .A2(n5151), .ZN(n5188) );
  NAND2_X2 U331 ( .A1(n4781), .A2(n33), .ZN(n4785) );
  INV_X2 U337 ( .A(n5260), .ZN(n454) );
  NAND2_X2 U339 ( .A1(n37), .A2(n5174), .ZN(n5252) );
  NAND2_X2 U340 ( .A1(n5173), .A2(n1042), .ZN(n37) );
  NAND2_X2 U341 ( .A1(n38), .A2(n2518), .ZN(n1088) );
  NAND2_X2 U342 ( .A1(n2826), .A2(n2410), .ZN(n2518) );
  NAND2_X2 U343 ( .A1(n6214), .A2(n1041), .ZN(n38) );
  NOR2_X2 U345 ( .A1(n5930), .A2(n259), .ZN(n6134) );
  NOR2_X4 U346 ( .A1(n5255), .A2(n5253), .ZN(n2291) );
  NOR2_X2 U347 ( .A1(n5171), .A2(n5172), .ZN(n5253) );
  INV_X4 U348 ( .A(n39), .ZN(n5255) );
  NAND2_X2 U349 ( .A1(n5171), .A2(n5172), .ZN(n39) );
  BUF_X4 U351 ( .A(n5295), .Z(n41) );
  NAND2_X2 U352 ( .A1(n6513), .A2(n4895), .ZN(n433) );
  OAI22_X2 U353 ( .A1(n1060), .A2(b[7]), .B1(n805), .B2(n2143), .ZN(n1980) );
  AOI22_X2 U356 ( .A1(n1107), .A2(n4614), .B1(n1194), .B2(b[13]), .ZN(n1191)
         );
  NAND2_X2 U360 ( .A1(n44), .A2(n661), .ZN(n2398) );
  NAND2_X2 U361 ( .A1(n659), .A2(n660), .ZN(n44) );
  NAND2_X2 U363 ( .A1(n4824), .A2(n1063), .ZN(n2371) );
  NOR2_X2 U364 ( .A1(n45), .A2(n5555), .ZN(n1724) );
  INV_X2 U365 ( .A(n5557), .ZN(n45) );
  NAND2_X2 U366 ( .A1(n2520), .A2(n2522), .ZN(n5557) );
  NAND2_X2 U368 ( .A1(n5094), .A2(n3466), .ZN(n2767) );
  NAND2_X1 U373 ( .A1(n6221), .A2(n1060), .ZN(n2644) );
  NAND2_X2 U378 ( .A1(n49), .A2(n2692), .ZN(n2694) );
  INV_X2 U379 ( .A(n2769), .ZN(n49) );
  NAND2_X2 U380 ( .A1(n562), .A2(n561), .ZN(n2769) );
  NAND2_X2 U381 ( .A1(n1996), .A2(n4650), .ZN(n1994) );
  NAND2_X2 U382 ( .A1(n2694), .A2(n2693), .ZN(n1846) );
  NAND2_X2 U384 ( .A1(n3126), .A2(n5804), .ZN(n3672) );
  AOI22_X2 U385 ( .A1(n1079), .A2(n1667), .B1(n3602), .B2(n3603), .ZN(n5804)
         );
  NAND2_X2 U386 ( .A1(n1081), .A2(n1080), .ZN(n3126) );
  NOR3_X4 U387 ( .A1(n50), .A2(n2767), .A3(n5320), .ZN(n5596) );
  NAND3_X2 U388 ( .A1(n5919), .A2(n628), .A3(n343), .ZN(n50) );
  NAND2_X2 U393 ( .A1(n1985), .A2(n1984), .ZN(n4912) );
  NAND2_X2 U394 ( .A1(n895), .A2(n894), .ZN(n1985) );
  INV_X4 U397 ( .A(n337), .ZN(n4071) );
  NAND2_X4 U398 ( .A1(n1295), .A2(n1294), .ZN(n337) );
  OAI21_X2 U399 ( .B1(n4759), .B2(n4758), .A(n2321), .ZN(n1788) );
  AOI22_X2 U402 ( .A1(n3869), .A2(a[0]), .B1(n4219), .B2(n984), .ZN(n3912) );
  NAND2_X2 U404 ( .A1(n3448), .A2(n3447), .ZN(n2374) );
  INV_X4 U405 ( .A(n51), .ZN(n3482) );
  NAND2_X2 U407 ( .A1(n2110), .A2(n2111), .ZN(n485) );
  NOR2_X2 U408 ( .A1(n3706), .A2(n3745), .ZN(n2111) );
  NAND3_X2 U409 ( .A1(n1458), .A2(n3521), .A3(n3523), .ZN(n3350) );
  NAND2_X2 U410 ( .A1(n1641), .A2(n3524), .ZN(n3521) );
  NAND2_X2 U411 ( .A1(n53), .A2(n6151), .ZN(n1338) );
  NAND2_X2 U413 ( .A1(n3491), .A2(n281), .ZN(n53) );
  NAND2_X2 U415 ( .A1(n2298), .A2(n3983), .ZN(n2238) );
  BUF_X4 U416 ( .A(n3304), .Z(n54) );
  NAND2_X2 U421 ( .A1(n55), .A2(n3289), .ZN(n194) );
  INV_X2 U422 ( .A(n2383), .ZN(n55) );
  NAND2_X2 U423 ( .A1(n697), .A2(n696), .ZN(n2383) );
  NOR2_X4 U425 ( .A1(a[11]), .A2(a[12]), .ZN(n2473) );
  NAND2_X2 U429 ( .A1(n6000), .A2(n5609), .ZN(n5616) );
  NOR2_X2 U430 ( .A1(n6200), .A2(n1943), .ZN(n172) );
  INV_X4 U432 ( .A(n4882), .ZN(n1440) );
  NOR2_X2 U436 ( .A1(n2583), .A2(n3474), .ZN(n3396) );
  NAND2_X2 U437 ( .A1(n699), .A2(n3538), .ZN(n1933) );
  NAND2_X2 U438 ( .A1(n337), .A2(n4073), .ZN(n819) );
  NAND2_X2 U442 ( .A1(n2500), .A2(n2849), .ZN(n3557) );
  NAND2_X2 U443 ( .A1(n3011), .A2(n5360), .ZN(n2502) );
  NAND2_X4 U444 ( .A1(n6654), .A2(a[13]), .ZN(n3011) );
  NAND2_X2 U446 ( .A1(n4692), .A2(n245), .ZN(n993) );
  NOR2_X2 U448 ( .A1(n4890), .A2(n59), .ZN(n4921) );
  NOR2_X2 U449 ( .A1(n5190), .A2(n4889), .ZN(n59) );
  NAND2_X2 U451 ( .A1(n1798), .A2(n1800), .ZN(n5019) );
  NAND2_X2 U453 ( .A1(n824), .A2(n823), .ZN(n1507) );
  BUF_X4 U454 ( .A(n2757), .Z(n60) );
  BUF_X4 U456 ( .A(n6086), .Z(n61) );
  NAND2_X2 U457 ( .A1(n3161), .A2(n3342), .ZN(n1102) );
  NAND2_X2 U458 ( .A1(n2326), .A2(n4558), .ZN(n1276) );
  NOR2_X2 U460 ( .A1(n4217), .A2(b[3]), .ZN(n1775) );
  NOR2_X2 U461 ( .A1(n1775), .A2(n1774), .ZN(n1773) );
  INV_X4 U462 ( .A(n4657), .ZN(n2546) );
  NAND3_X2 U463 ( .A1(n993), .A2(n3130), .A3(n3129), .ZN(n3127) );
  AOI22_X2 U465 ( .A1(n6450), .A2(n1457), .B1(n4529), .B2(n4408), .ZN(n2995)
         );
  NAND2_X2 U468 ( .A1(n4042), .A2(n4040), .ZN(n63) );
  OAI21_X2 U471 ( .B1(n3775), .B2(n3776), .A(n66), .ZN(n3778) );
  NAND2_X2 U472 ( .A1(n6161), .A2(n6445), .ZN(n66) );
  NAND2_X2 U475 ( .A1(n1911), .A2(n1910), .ZN(n1534) );
  OAI21_X2 U476 ( .B1(n1913), .B2(n1912), .A(n3654), .ZN(n1910) );
  BUF_X4 U477 ( .A(n5694), .Z(n69) );
  NAND2_X2 U479 ( .A1(n2508), .A2(n4231), .ZN(n70) );
  NAND3_X2 U480 ( .A1(n71), .A2(n4338), .A3(n2180), .ZN(n4488) );
  NAND2_X2 U481 ( .A1(n990), .A2(n2081), .ZN(n71) );
  INV_X4 U482 ( .A(n72), .ZN(n1140) );
  NOR2_X2 U483 ( .A1(n6186), .A2(n2602), .ZN(n72) );
  NAND2_X2 U484 ( .A1(n73), .A2(n349), .ZN(n4069) );
  NAND2_X2 U485 ( .A1(n347), .A2(n348), .ZN(n73) );
  INV_X4 U486 ( .A(n3617), .ZN(n3052) );
  NAND2_X2 U487 ( .A1(n4582), .A2(n2130), .ZN(n2167) );
  OAI22_X2 U489 ( .A1(n74), .A2(n4300), .B1(n4298), .B2(n1320), .ZN(n5717) );
  NOR2_X2 U490 ( .A1(n4296), .A2(n4297), .ZN(n74) );
  XOR2_X2 U492 ( .A(b[8]), .B(a[9]), .Z(n75) );
  INV_X4 U493 ( .A(n1914), .ZN(n1911) );
  NAND2_X2 U500 ( .A1(n78), .A2(n779), .ZN(n3073) );
  NAND2_X2 U501 ( .A1(n777), .A2(n4721), .ZN(n78) );
  NOR2_X2 U502 ( .A1(n4578), .A2(n4577), .ZN(n4580) );
  NAND2_X2 U504 ( .A1(n1759), .A2(n5212), .ZN(n823) );
  INV_X4 U508 ( .A(n4514), .ZN(n4517) );
  NOR2_X2 U509 ( .A1(n758), .A2(n2249), .ZN(n3175) );
  NAND3_X2 U510 ( .A1(n1448), .A2(a[19]), .A3(a[20]), .ZN(n758) );
  NOR2_X2 U511 ( .A1(n4356), .A2(n80), .ZN(n4404) );
  NAND2_X2 U512 ( .A1(n83), .A2(n81), .ZN(n80) );
  NAND2_X2 U513 ( .A1(n1194), .A2(b[4]), .ZN(n81) );
  NAND2_X2 U515 ( .A1(n1193), .A2(n4598), .ZN(n83) );
  NAND3_X2 U516 ( .A1(n3308), .A2(a[19]), .A3(n5471), .ZN(n5364) );
  NAND3_X2 U518 ( .A1(n3285), .A2(n1976), .A3(n3078), .ZN(n84) );
  INV_X2 U523 ( .A(n5718), .ZN(n2235) );
  INV_X4 U524 ( .A(n86), .ZN(n1753) );
  NOR2_X2 U525 ( .A1(n1754), .A2(n4479), .ZN(n86) );
  INV_X4 U526 ( .A(n4584), .ZN(n1997) );
  XNOR2_X2 U528 ( .A(n3650), .B(n3901), .ZN(n2649) );
  NAND2_X2 U529 ( .A1(n4637), .A2(n4635), .ZN(n2226) );
  XNOR2_X2 U530 ( .A(n1110), .B(n4476), .ZN(n4637) );
  NAND2_X1 U533 ( .A1(n998), .A2(n4614), .ZN(n87) );
  NAND2_X2 U534 ( .A1(n757), .A2(n756), .ZN(n3064) );
  NAND3_X2 U535 ( .A1(n2081), .A2(n88), .A3(n2090), .ZN(n1157) );
  NOR2_X2 U537 ( .A1(n3731), .A2(n2131), .ZN(n2092) );
  INV_X2 U538 ( .A(n2324), .ZN(n754) );
  NAND2_X2 U539 ( .A1(n279), .A2(n278), .ZN(n2324) );
  NAND2_X2 U540 ( .A1(n89), .A2(n4005), .ZN(n697) );
  INV_X2 U541 ( .A(n4293), .ZN(n89) );
  AOI21_X2 U546 ( .B1(n3941), .B2(n6558), .A(n91), .ZN(n4056) );
  NAND2_X2 U547 ( .A1(n94), .A2(n92), .ZN(n91) );
  NAND2_X2 U550 ( .A1(n4506), .A2(b[13]), .ZN(n94) );
  NAND2_X2 U551 ( .A1(n95), .A2(n791), .ZN(n793) );
  INV_X2 U552 ( .A(n3974), .ZN(n95) );
  NOR3_X2 U553 ( .A1(n992), .A2(n988), .A3(n3904), .ZN(n3974) );
  INV_X4 U554 ( .A(n4376), .ZN(n2347) );
  NAND3_X1 U555 ( .A1(n690), .A2(n432), .A3(n2929), .ZN(n931) );
  NAND2_X2 U556 ( .A1(n4515), .A2(n4512), .ZN(n2325) );
  INV_X4 U560 ( .A(n4612), .ZN(n3568) );
  INV_X4 U562 ( .A(n96), .ZN(n1848) );
  NOR2_X4 U563 ( .A1(n2469), .A2(n1417), .ZN(n96) );
  NAND2_X2 U564 ( .A1(n525), .A2(n524), .ZN(n1077) );
  NAND2_X2 U569 ( .A1(n98), .A2(n2243), .ZN(n1079) );
  NAND2_X2 U572 ( .A1(n319), .A2(n3409), .ZN(n930) );
  NOR2_X2 U576 ( .A1(n101), .A2(n100), .ZN(n2818) );
  NOR2_X2 U577 ( .A1(n2491), .A2(n254), .ZN(n100) );
  NOR2_X2 U578 ( .A1(n4670), .A2(n54), .ZN(n101) );
  NAND2_X2 U579 ( .A1(n2156), .A2(n1098), .ZN(n2152) );
  OAI21_X2 U580 ( .B1(n1710), .B2(n2042), .A(n3331), .ZN(n2646) );
  NAND2_X2 U581 ( .A1(n4563), .A2(n4564), .ZN(n444) );
  OAI21_X2 U583 ( .B1(n1006), .B2(n3408), .A(n2803), .ZN(n1582) );
  AOI21_X2 U584 ( .B1(n1004), .B2(n4486), .A(n3051), .ZN(n2803) );
  INV_X4 U585 ( .A(n4576), .ZN(n1006) );
  INV_X4 U588 ( .A(n4564), .ZN(n442) );
  NAND2_X2 U590 ( .A1(n2411), .A2(n6402), .ZN(n676) );
  NAND2_X2 U592 ( .A1(n677), .A2(n676), .ZN(n5324) );
  XNOR2_X2 U593 ( .A(n103), .B(n5027), .ZN(n2757) );
  AOI22_X2 U594 ( .A1(n6452), .A2(n2750), .B1(n1619), .B2(n1035), .ZN(n103) );
  INV_X4 U595 ( .A(n4563), .ZN(n443) );
  NOR2_X2 U596 ( .A1(n6022), .A2(n1145), .ZN(n6023) );
  NAND3_X2 U597 ( .A1(n1781), .A2(n1780), .A3(n5111), .ZN(n1779) );
  NOR2_X2 U600 ( .A1(n6569), .A2(n4601), .ZN(n3664) );
  NAND2_X2 U601 ( .A1(n1506), .A2(n5210), .ZN(n509) );
  NAND2_X2 U602 ( .A1(n3308), .A2(n2749), .ZN(n3624) );
  NAND2_X2 U603 ( .A1(n4689), .A2(b[21]), .ZN(n4816) );
  NAND2_X4 U604 ( .A1(a[23]), .A2(b[6]), .ZN(n4924) );
  NAND2_X2 U609 ( .A1(n611), .A2(n585), .ZN(n2272) );
  NAND2_X2 U610 ( .A1(n108), .A2(n5032), .ZN(n5038) );
  NAND2_X2 U611 ( .A1(n2600), .A2(n2599), .ZN(n108) );
  NAND2_X2 U612 ( .A1(n1540), .A2(n1685), .ZN(n875) );
  INV_X2 U614 ( .A(n2063), .ZN(n1721) );
  NAND2_X2 U615 ( .A1(n2064), .A2(n2810), .ZN(n2063) );
  NOR2_X2 U618 ( .A1(n5930), .A2(n5929), .ZN(n2330) );
  NAND3_X2 U619 ( .A1(n5926), .A2(n6005), .A3(n1675), .ZN(n5930) );
  NAND2_X4 U620 ( .A1(n916), .A2(n1024), .ZN(n2218) );
  NAND2_X4 U622 ( .A1(n809), .A2(n810), .ZN(n812) );
  NAND2_X2 U623 ( .A1(n111), .A2(n110), .ZN(n1907) );
  NAND2_X2 U624 ( .A1(n1941), .A2(n5039), .ZN(n110) );
  NAND2_X2 U625 ( .A1(n1112), .A2(n1942), .ZN(n111) );
  NOR2_X4 U626 ( .A1(n5190), .A2(n4604), .ZN(n3085) );
  NAND2_X2 U628 ( .A1(n4481), .A2(n1127), .ZN(n1930) );
  NAND2_X2 U630 ( .A1(n116), .A2(n114), .ZN(n113) );
  NAND2_X2 U631 ( .A1(n2406), .A2(b[19]), .ZN(n114) );
  NOR2_X2 U636 ( .A1(n1992), .A2(n1991), .ZN(n4734) );
  NAND2_X2 U640 ( .A1(n117), .A2(n1380), .ZN(n1336) );
  NAND2_X2 U641 ( .A1(n418), .A2(n419), .ZN(n117) );
  NAND2_X2 U643 ( .A1(n1193), .A2(n5277), .ZN(n118) );
  NAND2_X2 U647 ( .A1(n737), .A2(n738), .ZN(n119) );
  NAND2_X2 U649 ( .A1(n3500), .A2(n646), .ZN(n120) );
  NAND2_X2 U655 ( .A1(n4488), .A2(n787), .ZN(n2530) );
  NOR2_X2 U658 ( .A1(n2331), .A2(n2330), .ZN(n388) );
  NAND2_X2 U662 ( .A1(n123), .A2(n4528), .ZN(n1600) );
  NAND2_X2 U663 ( .A1(n2691), .A2(n2690), .ZN(n123) );
  NAND2_X2 U664 ( .A1(n3832), .A2(n2276), .ZN(n2275) );
  OAI21_X2 U665 ( .B1(n1957), .B2(n124), .A(n4838), .ZN(n1224) );
  NAND2_X2 U667 ( .A1(n4839), .A2(n1226), .ZN(n2348) );
  NAND2_X2 U670 ( .A1(n2051), .A2(n2050), .ZN(n125) );
  INV_X2 U673 ( .A(n1270), .ZN(n127) );
  NAND3_X1 U675 ( .A1(n3670), .A2(n5862), .A3(n2879), .ZN(n5867) );
  NOR2_X4 U676 ( .A1(n5314), .A2(n3105), .ZN(n3670) );
  NAND2_X2 U678 ( .A1(n2044), .A2(n5069), .ZN(n3524) );
  INV_X4 U687 ( .A(n2468), .ZN(n1285) );
  NAND2_X2 U688 ( .A1(n132), .A2(n2189), .ZN(n2295) );
  NAND2_X2 U689 ( .A1(n3937), .A2(n3938), .ZN(n132) );
  OAI21_X2 U691 ( .B1(n280), .B2(n2517), .A(n5133), .ZN(n133) );
  NAND2_X2 U692 ( .A1(n2468), .A2(n5014), .ZN(n5069) );
  NAND2_X2 U693 ( .A1(n136), .A2(n134), .ZN(n5058) );
  NAND2_X2 U696 ( .A1(n6035), .A2(n865), .ZN(n136) );
  NAND2_X2 U699 ( .A1(n137), .A2(n691), .ZN(n1716) );
  NAND2_X2 U700 ( .A1(n689), .A2(n690), .ZN(n137) );
  OAI21_X2 U701 ( .B1(n1714), .B2(n1530), .A(n6391), .ZN(n1713) );
  NAND2_X2 U702 ( .A1(n1240), .A2(n4901), .ZN(n2219) );
  NAND2_X2 U703 ( .A1(n595), .A2(n594), .ZN(n4901) );
  NAND3_X1 U704 ( .A1(n256), .A2(n6525), .A3(n3758), .ZN(n5593) );
  BUF_X4 U710 ( .A(n4805), .Z(n139) );
  NOR2_X2 U712 ( .A1(n2936), .A2(n5389), .ZN(n5388) );
  NAND2_X4 U713 ( .A1(n1164), .A2(n1163), .ZN(n4760) );
  NAND2_X2 U714 ( .A1(n2143), .A2(n328), .ZN(n1091) );
  NAND2_X2 U716 ( .A1(n141), .A2(n140), .ZN(n3275) );
  NAND2_X2 U719 ( .A1(n142), .A2(n1321), .ZN(n1925) );
  BUF_X4 U721 ( .A(n5729), .Z(n143) );
  NAND2_X2 U723 ( .A1(n1753), .A2(n1752), .ZN(n1594) );
  NAND2_X2 U726 ( .A1(n4589), .A2(n1529), .ZN(n2470) );
  NAND2_X2 U729 ( .A1(n3727), .A2(n4720), .ZN(n1437) );
  NAND2_X2 U730 ( .A1(n4656), .A2(n4655), .ZN(n3727) );
  NOR3_X2 U731 ( .A1(n1339), .A2(n5886), .A3(n145), .ZN(\d[42]_BAR ) );
  NOR3_X1 U732 ( .A1(n6062), .A2(n5876), .A3(n5884), .ZN(n145) );
  BUF_X4 U733 ( .A(n4736), .Z(n146) );
  OAI21_X2 U734 ( .B1(n3073), .B2(n146), .A(n1350), .ZN(n1376) );
  NOR2_X2 U735 ( .A1(n4975), .A2(n2949), .ZN(n5839) );
  INV_X4 U736 ( .A(n2975), .ZN(n2974) );
  NAND2_X2 U737 ( .A1(n4762), .A2(n4760), .ZN(n3129) );
  INV_X2 U740 ( .A(n4917), .ZN(n573) );
  NAND2_X2 U741 ( .A1(n1376), .A2(n1375), .ZN(n4917) );
  INV_X4 U743 ( .A(n2488), .ZN(n1653) );
  NAND2_X2 U746 ( .A1(n3253), .A2(n3713), .ZN(n148) );
  OAI21_X2 U747 ( .B1(n1653), .B2(n2384), .A(n1844), .ZN(n2469) );
  NAND2_X4 U748 ( .A1(n150), .A2(n149), .ZN(n1844) );
  INV_X4 U749 ( .A(n1845), .ZN(n149) );
  INV_X4 U750 ( .A(n1846), .ZN(n150) );
  OAI22_X2 U752 ( .A1(n1683), .A2(n4904), .B1(n4906), .B2(n4905), .ZN(n1984)
         );
  AOI22_X2 U755 ( .A1(n3074), .A2(n3077), .B1(n5039), .B2(n6202), .ZN(n3273)
         );
  NOR2_X4 U756 ( .A1(n1461), .A2(n5099), .ZN(n5377) );
  NOR2_X2 U761 ( .A1(n154), .A2(n2630), .ZN(n3247) );
  NOR2_X2 U767 ( .A1(n2700), .A2(n3080), .ZN(n4539) );
  NAND2_X2 U769 ( .A1(n6377), .A2(n2852), .ZN(n1947) );
  NAND2_X2 U771 ( .A1(n3157), .A2(n6059), .ZN(n6055) );
  NAND2_X4 U773 ( .A1(n2219), .A2(n2218), .ZN(n3074) );
  INV_X1 U774 ( .A(n3726), .ZN(n2278) );
  INV_X4 U775 ( .A(n3645), .ZN(n4655) );
  NAND2_X2 U777 ( .A1(n4599), .A2(n586), .ZN(n1546) );
  NAND2_X4 U779 ( .A1(n1202), .A2(n162), .ZN(n1417) );
  NAND2_X2 U780 ( .A1(n1850), .A2(n1465), .ZN(n162) );
  BUF_X4 U781 ( .A(n5647), .Z(n163) );
  NOR2_X2 U782 ( .A1(n3113), .A2(n3114), .ZN(n1500) );
  NAND2_X2 U783 ( .A1(n1502), .A2(n1501), .ZN(n3113) );
  NOR2_X4 U784 ( .A1(n217), .A2(b[14]), .ZN(n4592) );
  NAND3_X2 U785 ( .A1(n2313), .A2(n2314), .A3(n2315), .ZN(n4833) );
  NAND2_X2 U786 ( .A1(n3385), .A2(n3469), .ZN(n2313) );
  NAND2_X2 U790 ( .A1(n2643), .A2(n2642), .ZN(n164) );
  NAND4_X1 U791 ( .A1(n165), .A2(n5392), .A3(n5393), .A4(n5391), .ZN(
        \d[33]_BAR ) );
  NAND3_X2 U792 ( .A1(n1327), .A2(n345), .A3(n5390), .ZN(n165) );
  NOR2_X2 U794 ( .A1(n3724), .A2(n3359), .ZN(n4982) );
  AOI22_X2 U795 ( .A1(n4409), .A2(n564), .B1(n4410), .B2(n4411), .ZN(n4412) );
  NOR2_X2 U796 ( .A1(n4070), .A2(n818), .ZN(n2973) );
  AOI22_X2 U797 ( .A1(n5360), .A2(n2510), .B1(n2382), .B2(b[18]), .ZN(n5169)
         );
  NOR2_X2 U799 ( .A1(n5034), .A2(n166), .ZN(n2597) );
  NAND2_X2 U800 ( .A1(n3090), .A2(n3089), .ZN(n166) );
  INV_X4 U801 ( .A(n5458), .ZN(n1344) );
  NAND2_X2 U803 ( .A1(n4895), .A2(n6513), .ZN(n167) );
  NAND3_X2 U804 ( .A1(n6000), .A2(n5995), .A3(n6068), .ZN(n5931) );
  NAND2_X2 U808 ( .A1(n5508), .A2(n972), .ZN(n2069) );
  NAND2_X2 U809 ( .A1(n169), .A2(n168), .ZN(n972) );
  INV_X2 U810 ( .A(n5553), .ZN(n168) );
  INV_X2 U811 ( .A(n5552), .ZN(n169) );
  NAND2_X2 U812 ( .A1(n1267), .A2(n1265), .ZN(n3155) );
  AOI22_X2 U813 ( .A1(n1778), .A2(n952), .B1(n538), .B2(n780), .ZN(n1267) );
  NAND2_X2 U817 ( .A1(n214), .A2(n2403), .ZN(n4338) );
  AOI21_X2 U822 ( .B1(n1769), .B2(n4650), .A(n4651), .ZN(n4735) );
  NAND2_X2 U823 ( .A1(n4520), .A2(n4519), .ZN(n4573) );
  NAND2_X2 U827 ( .A1(n192), .A2(n1504), .ZN(n3114) );
  NAND2_X2 U831 ( .A1(n1176), .A2(n173), .ZN(n3986) );
  NAND2_X1 U832 ( .A1(n1175), .A2(n3984), .ZN(n173) );
  NAND2_X2 U833 ( .A1(n4277), .A2(n4279), .ZN(n2208) );
  NAND2_X2 U834 ( .A1(n3843), .A2(n3842), .ZN(n4277) );
  NAND2_X2 U836 ( .A1(n3009), .A2(n1257), .ZN(n3008) );
  NAND2_X2 U837 ( .A1(n2508), .A2(n4231), .ZN(n1149) );
  NAND2_X4 U838 ( .A1(n1140), .A2(n2506), .ZN(n2508) );
  NAND2_X2 U839 ( .A1(n939), .A2(n940), .ZN(n174) );
  NOR2_X2 U840 ( .A1(n3076), .A2(n6587), .ZN(n2847) );
  NAND2_X2 U841 ( .A1(n1013), .A2(n5984), .ZN(n5973) );
  NAND2_X2 U842 ( .A1(n657), .A2(n658), .ZN(n4158) );
  NAND2_X2 U843 ( .A1(n175), .A2(n4247), .ZN(n4285) );
  NAND3_X2 U844 ( .A1(n1551), .A2(n1553), .A3(n4245), .ZN(n175) );
  INV_X2 U845 ( .A(n2172), .ZN(n268) );
  NAND2_X2 U846 ( .A1(n620), .A2(n619), .ZN(n2172) );
  INV_X2 U847 ( .A(n5305), .ZN(n176) );
  AOI21_X2 U848 ( .B1(n5303), .B2(n5302), .A(n5301), .ZN(n5305) );
  NAND2_X1 U849 ( .A1(n3286), .A2(n4295), .ZN(n2831) );
  NAND2_X2 U850 ( .A1(n2669), .A2(n2668), .ZN(n4295) );
  NAND2_X2 U851 ( .A1(n2964), .A2(n2321), .ZN(n2963) );
  INV_X4 U852 ( .A(n177), .ZN(n339) );
  XNOR2_X2 U855 ( .A(n178), .B(n5457), .ZN(n2522) );
  NAND2_X2 U856 ( .A1(n387), .A2(n386), .ZN(n178) );
  NAND2_X2 U857 ( .A1(n548), .A2(n179), .ZN(n550) );
  XNOR2_X2 U859 ( .A(n2971), .B(n1008), .ZN(n1136) );
  NAND2_X2 U863 ( .A1(n1355), .A2(n5975), .ZN(n5970) );
  NAND2_X2 U865 ( .A1(n2099), .A2(n3024), .ZN(n448) );
  NOR2_X2 U867 ( .A1(n5143), .A2(n5056), .ZN(n181) );
  AOI21_X2 U870 ( .B1(n4194), .B2(n4193), .A(n4192), .ZN(n5689) );
  NAND2_X2 U871 ( .A1(n183), .A2(n182), .ZN(n5139) );
  NAND2_X2 U872 ( .A1(n5136), .A2(b[13]), .ZN(n182) );
  OR2_X2 U876 ( .A1(n1847), .A2(b[2]), .ZN(n2248) );
  INV_X4 U879 ( .A(n1969), .ZN(n1038) );
  NAND2_X2 U880 ( .A1(n2383), .A2(n4295), .ZN(n911) );
  INV_X2 U881 ( .A(n3211), .ZN(n857) );
  NAND2_X2 U886 ( .A1(n699), .A2(n6569), .ZN(n3591) );
  NAND2_X2 U887 ( .A1(n4307), .A2(n2242), .ZN(n2241) );
  INV_X2 U888 ( .A(n4267), .ZN(n3364) );
  NAND2_X2 U890 ( .A1(n2173), .A2(n4300), .ZN(n842) );
  NAND2_X2 U893 ( .A1(n4229), .A2(n4228), .ZN(n1123) );
  NAND2_X2 U896 ( .A1(n3588), .A2(n3589), .ZN(n2388) );
  NAND2_X2 U897 ( .A1(n3213), .A2(n2389), .ZN(n3588) );
  NAND2_X2 U899 ( .A1(n1200), .A2(n1197), .ZN(n4667) );
  NAND2_X2 U901 ( .A1(n1279), .A2(n1280), .ZN(n2179) );
  INV_X2 U907 ( .A(n2511), .ZN(n190) );
  INV_X2 U913 ( .A(n4470), .ZN(n2366) );
  AOI21_X2 U914 ( .B1(n3853), .B2(n6558), .A(n3852), .ZN(n3892) );
  NAND2_X2 U916 ( .A1(n1159), .A2(n1158), .ZN(n3303) );
  BUF_X4 U919 ( .A(n6035), .Z(n195) );
  INV_X2 U920 ( .A(n1873), .ZN(n1370) );
  NAND2_X2 U921 ( .A1(n601), .A2(n3095), .ZN(n1873) );
  XNOR2_X2 U923 ( .A(n3087), .B(n4469), .ZN(n1842) );
  NAND2_X2 U925 ( .A1(n196), .A2(n731), .ZN(n3192) );
  NAND2_X2 U926 ( .A1(n729), .A2(n5558), .ZN(n196) );
  NAND2_X2 U928 ( .A1(n5924), .A2(n3389), .ZN(n4977) );
  NAND2_X2 U929 ( .A1(n197), .A2(n2458), .ZN(n2457) );
  NOR2_X2 U930 ( .A1(n2460), .A2(n2467), .ZN(n197) );
  NAND2_X2 U931 ( .A1(n3457), .A2(n4183), .ZN(n3456) );
  NAND2_X2 U932 ( .A1(n199), .A2(n198), .ZN(n4185) );
  NAND2_X2 U934 ( .A1(n4506), .A2(b[4]), .ZN(n199) );
  NAND2_X2 U936 ( .A1(n202), .A2(n201), .ZN(n4353) );
  NAND2_X2 U938 ( .A1(n1127), .A2(n4346), .ZN(n202) );
  NOR2_X4 U940 ( .A1(n1603), .A2(a[19]), .ZN(n5894) );
  INV_X8 U941 ( .A(a[21]), .ZN(n1603) );
  XNOR2_X2 U942 ( .A(n5554), .B(n5553), .ZN(n5562) );
  OAI21_X1 U943 ( .B1(n4995), .B2(b[3]), .A(n6158), .ZN(n4401) );
  NAND2_X2 U946 ( .A1(n1147), .A2(b[3]), .ZN(n1932) );
  INV_X4 U947 ( .A(n4794), .ZN(n4810) );
  OAI21_X2 U950 ( .B1(n206), .B2(n5055), .A(n1515), .ZN(n5143) );
  AOI22_X2 U951 ( .A1(n1516), .A2(n1517), .B1(n282), .B2(n5053), .ZN(n206) );
  NOR2_X2 U954 ( .A1(n1749), .A2(n1748), .ZN(n1747) );
  NAND2_X2 U955 ( .A1(n1639), .A2(n1638), .ZN(n3523) );
  NAND2_X2 U956 ( .A1(n5049), .A2(n5047), .ZN(n5045) );
  NAND2_X2 U957 ( .A1(n5042), .A2(n5044), .ZN(n5047) );
  NAND2_X2 U960 ( .A1(n510), .A2(n509), .ZN(n1627) );
  AOI22_X2 U961 ( .A1(n4409), .A2(n564), .B1(n4410), .B2(n4411), .ZN(n327) );
  NAND3_X2 U962 ( .A1(n208), .A2(n1962), .A3(n4075), .ZN(n1961) );
  INV_X2 U963 ( .A(n3980), .ZN(n208) );
  OAI21_X2 U964 ( .B1(n2973), .B2(n4071), .A(n2972), .ZN(n3980) );
  NOR3_X2 U965 ( .A1(n6017), .A2(n5381), .A3(n6205), .ZN(n6021) );
  INV_X4 U966 ( .A(b[23]), .ZN(n979) );
  NAND2_X2 U967 ( .A1(n1974), .A2(n5091), .ZN(n2421) );
  NOR2_X4 U969 ( .A1(a[5]), .A2(a[6]), .ZN(n3877) );
  NAND2_X2 U971 ( .A1(n3975), .A2(n3974), .ZN(n792) );
  AOI21_X2 U973 ( .B1(n978), .B2(a[9]), .A(n3636), .ZN(n3635) );
  NAND2_X2 U975 ( .A1(n5144), .A2(n2108), .ZN(n5056) );
  NAND2_X4 U977 ( .A1(n3991), .A2(a[11]), .ZN(n998) );
  NAND2_X2 U981 ( .A1(n211), .A2(n210), .ZN(n2005) );
  NAND2_X2 U983 ( .A1(n788), .A2(n789), .ZN(n211) );
  INV_X4 U986 ( .A(n4486), .ZN(n4484) );
  NAND2_X2 U987 ( .A1(n1468), .A2(n1467), .ZN(n664) );
  NAND2_X4 U988 ( .A1(n213), .A2(n702), .ZN(n4776) );
  NAND2_X4 U989 ( .A1(n700), .A2(n701), .ZN(n213) );
  NAND2_X2 U992 ( .A1(n892), .A2(n4869), .ZN(n895) );
  NAND2_X2 U996 ( .A1(n2182), .A2(n2181), .ZN(n214) );
  NAND2_X2 U997 ( .A1(n215), .A2(n1027), .ZN(n2163) );
  NAND2_X1 U998 ( .A1(n2083), .A2(n3580), .ZN(n215) );
  NOR2_X4 U1003 ( .A1(n2117), .A2(n3264), .ZN(n216) );
  INV_X4 U1004 ( .A(n998), .ZN(n217) );
  NOR2_X2 U1005 ( .A1(n217), .A2(b[3]), .ZN(n3775) );
  NOR2_X2 U1006 ( .A1(n3778), .A2(n1225), .ZN(n1511) );
  NAND2_X2 U1009 ( .A1(n2166), .A2(n2479), .ZN(n2601) );
  AOI21_X2 U1013 ( .B1(n3086), .B2(n4545), .A(n3085), .ZN(n4624) );
  NAND2_X2 U1014 ( .A1(n218), .A2(n655), .ZN(n3283) );
  NAND2_X2 U1015 ( .A1(n653), .A2(n654), .ZN(n218) );
  NOR2_X4 U1016 ( .A1(n1612), .A2(n5489), .ZN(n1610) );
  NAND2_X2 U1018 ( .A1(n758), .A2(b[4]), .ZN(n2540) );
  NOR2_X2 U1021 ( .A1(n5451), .A2(n5450), .ZN(n5452) );
  NAND2_X2 U1022 ( .A1(n5553), .A2(n5506), .ZN(n1179) );
  NAND2_X2 U1023 ( .A1(n221), .A2(n219), .ZN(n5276) );
  NAND2_X2 U1026 ( .A1(n309), .A2(b[21]), .ZN(n221) );
  NAND2_X2 U1027 ( .A1(n223), .A2(n222), .ZN(n5342) );
  NAND2_X2 U1028 ( .A1(n4767), .A2(n566), .ZN(n222) );
  NAND2_X4 U1031 ( .A1(n2435), .A2(n2434), .ZN(n2524) );
  NAND2_X4 U1032 ( .A1(n2032), .A2(a[20]), .ZN(n2435) );
  NAND2_X2 U1033 ( .A1(n998), .A2(n3263), .ZN(n3481) );
  INV_X4 U1036 ( .A(n2926), .ZN(n2917) );
  NAND2_X2 U1037 ( .A1(n2426), .A2(n3350), .ZN(n1974) );
  INV_X2 U1038 ( .A(n2130), .ZN(n1599) );
  NOR2_X4 U1044 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  INV_X4 U1045 ( .A(n5369), .ZN(n2812) );
  INV_X4 U1046 ( .A(n2072), .ZN(n5546) );
  NAND2_X2 U1048 ( .A1(n621), .A2(n622), .ZN(n228) );
  NAND2_X2 U1050 ( .A1(n652), .A2(n651), .ZN(n3083) );
  INV_X4 U1053 ( .A(n4365), .ZN(n4012) );
  NOR2_X2 U1055 ( .A1(n6214), .A2(n1041), .ZN(n229) );
  OAI22_X2 U1056 ( .A1(n1988), .A2(a[5]), .B1(n4740), .B2(n4821), .ZN(n3469)
         );
  OAI21_X2 U1060 ( .B1(n4668), .B2(n232), .A(n3221), .ZN(n2969) );
  NAND3_X1 U1063 ( .A1(n3407), .A2(n3551), .A3(n3389), .ZN(n3388) );
  NOR3_X2 U1064 ( .A1(n1274), .A2(n3552), .A3(n3553), .ZN(n3551) );
  OAI22_X2 U1066 ( .A1(n2309), .A2(n3872), .B1(n253), .B2(n3871), .ZN(n3911)
         );
  NAND2_X2 U1067 ( .A1(n234), .A2(n1833), .ZN(n1832) );
  NAND2_X2 U1068 ( .A1(n1835), .A2(n1834), .ZN(n234) );
  NAND2_X2 U1069 ( .A1(n235), .A2(n2461), .ZN(n1665) );
  NAND2_X2 U1070 ( .A1(n1022), .A2(n2837), .ZN(n235) );
  INV_X4 U1072 ( .A(n1267), .ZN(n1266) );
  NAND2_X2 U1073 ( .A1(n236), .A2(n852), .ZN(n5764) );
  NAND2_X2 U1074 ( .A1(n850), .A2(n851), .ZN(n236) );
  INV_X2 U1075 ( .A(n4474), .ZN(n534) );
  NAND2_X2 U1078 ( .A1(n3417), .A2(n3418), .ZN(n3420) );
  NAND3_X2 U1079 ( .A1(n238), .A2(n1185), .A3(n6446), .ZN(n3571) );
  NAND2_X2 U1083 ( .A1(n2347), .A2(n265), .ZN(n239) );
  NAND2_X4 U1088 ( .A1(n6614), .A2(a[13]), .ZN(n699) );
  NAND2_X2 U1089 ( .A1(n5326), .A2(n1016), .ZN(n2157) );
  AOI22_X2 U1090 ( .A1(n2086), .A2(n5834), .B1(n4641), .B2(n4640), .ZN(n5326)
         );
  NAND2_X2 U1091 ( .A1(n243), .A2(n241), .ZN(n5361) );
  NAND2_X1 U1092 ( .A1(n4829), .A2(b[17]), .ZN(n241) );
  NAND2_X2 U1094 ( .A1(n5526), .A2(n1212), .ZN(n243) );
  NOR2_X2 U1095 ( .A1(n5076), .A2(b[8]), .ZN(n4502) );
  NAND2_X2 U1097 ( .A1(n745), .A2(n744), .ZN(n244) );
  NOR2_X2 U1098 ( .A1(n5566), .A2(n5564), .ZN(n1723) );
  NAND2_X2 U1100 ( .A1(n3215), .A2(n4550), .ZN(n1882) );
  INV_X8 U1101 ( .A(a[2]), .ZN(n4674) );
  NAND2_X2 U1102 ( .A1(n4130), .A2(n246), .ZN(n4135) );
  NOR2_X2 U1103 ( .A1(n249), .A2(n247), .ZN(n246) );
  NOR2_X2 U1104 ( .A1(n4216), .A2(n248), .ZN(n247) );
  INV_X2 U1105 ( .A(b[1]), .ZN(n248) );
  NOR2_X2 U1106 ( .A1(n4217), .A2(b[1]), .ZN(n249) );
  XNOR2_X2 U1111 ( .A(a[10]), .B(a[9]), .ZN(n253) );
  INV_X1 U1114 ( .A(n1009), .ZN(n254) );
  OAI21_X2 U1118 ( .B1(n2952), .B2(n4316), .A(n260), .ZN(n5322) );
  INV_X1 U1119 ( .A(n4316), .ZN(n851) );
  NAND2_X2 U1120 ( .A1(n5526), .A2(n1324), .ZN(n2526) );
  NAND2_X2 U1122 ( .A1(n3208), .A2(n3209), .ZN(n255) );
  NAND2_X2 U1123 ( .A1(n3208), .A2(n3209), .ZN(n4549) );
  NAND2_X2 U1124 ( .A1(n5105), .A2(n4219), .ZN(n3208) );
  INV_X4 U1127 ( .A(n4526), .ZN(n257) );
  NAND2_X2 U1128 ( .A1(n827), .A2(n828), .ZN(n258) );
  NAND2_X2 U1131 ( .A1(n1909), .A2(n4315), .ZN(n260) );
  NAND2_X1 U1132 ( .A1(n2334), .A2(n2721), .ZN(n263) );
  NAND2_X2 U1133 ( .A1(n263), .A2(n264), .ZN(n3855) );
  NAND2_X1 U1136 ( .A1(n1909), .A2(n4315), .ZN(n2707) );
  INV_X4 U1137 ( .A(n4007), .ZN(n1909) );
  NAND2_X2 U1140 ( .A1(n712), .A2(n2223), .ZN(n265) );
  NAND2_X2 U1141 ( .A1(n712), .A2(n2223), .ZN(n4375) );
  INV_X1 U1142 ( .A(n4837), .ZN(n2834) );
  NAND2_X2 U1144 ( .A1(n2956), .A2(n4686), .ZN(n1509) );
  OAI21_X2 U1145 ( .B1(n3900), .B2(n3901), .A(n3650), .ZN(n266) );
  OAI21_X1 U1146 ( .B1(n3900), .B2(n3901), .A(n3650), .ZN(n3903) );
  NAND2_X1 U1148 ( .A1(n2172), .A2(n3554), .ZN(n270) );
  NAND2_X1 U1153 ( .A1(n5056), .A2(n5143), .ZN(n272) );
  NAND2_X2 U1155 ( .A1(n662), .A2(n663), .ZN(n665) );
  NAND2_X2 U1156 ( .A1(n6206), .A2(n4972), .ZN(n274) );
  NAND2_X2 U1157 ( .A1(n1343), .A2(n2107), .ZN(n275) );
  NAND2_X1 U1158 ( .A1(n2325), .A2(n4514), .ZN(n278) );
  NAND2_X2 U1159 ( .A1(n276), .A2(n4517), .ZN(n279) );
  INV_X2 U1160 ( .A(n2325), .ZN(n276) );
  NAND2_X2 U1162 ( .A1(n2107), .A2(n1343), .ZN(n3265) );
  INV_X4 U1164 ( .A(n430), .ZN(n2337) );
  NAND2_X4 U1165 ( .A1(n5996), .A2(n5995), .ZN(n6070) );
  NAND2_X2 U1167 ( .A1(n4551), .A2(n4552), .ZN(n281) );
  NAND2_X2 U1168 ( .A1(n4552), .A2(n4551), .ZN(n4669) );
  NOR2_X2 U1169 ( .A1(n2513), .A2(b[4]), .ZN(n4754) );
  INV_X8 U1170 ( .A(n5190), .ZN(n5010) );
  NAND2_X4 U1172 ( .A1(n3656), .A2(n3705), .ZN(n3453) );
  AOI21_X1 U1173 ( .B1(n4212), .B2(n4746), .A(b[0]), .ZN(n4214) );
  NAND2_X2 U1177 ( .A1(n2770), .A2(n808), .ZN(n5014) );
  NAND2_X1 U1181 ( .A1(n2550), .A2(n4248), .ZN(n288) );
  NOR2_X2 U1184 ( .A1(n1865), .A2(n4001), .ZN(n3811) );
  AOI21_X2 U1186 ( .B1(n3809), .B2(a[0]), .A(n3555), .ZN(n4001) );
  OAI21_X2 U1188 ( .B1(n1964), .B2(n4077), .A(n3980), .ZN(n1963) );
  NAND2_X2 U1190 ( .A1(n971), .A2(n1408), .ZN(n1412) );
  NOR2_X2 U1191 ( .A1(n2783), .A2(n2784), .ZN(n2779) );
  NAND2_X2 U1192 ( .A1(n2249), .A2(n328), .ZN(n4350) );
  NAND2_X2 U1193 ( .A1(n1868), .A2(n5789), .ZN(n290) );
  INV_X4 U1198 ( .A(n4605), .ZN(n1218) );
  NOR2_X2 U1199 ( .A1(n4605), .A2(n4604), .ZN(n4608) );
  XNOR2_X2 U1201 ( .A(n3860), .B(n3861), .ZN(n3024) );
  INV_X4 U1203 ( .A(n4913), .ZN(n419) );
  XOR2_X2 U1206 ( .A(a[3]), .B(b[19]), .Z(n2731) );
  NAND2_X1 U1207 ( .A1(n4322), .A2(n4323), .ZN(n293) );
  NOR2_X4 U1213 ( .A1(n3756), .A2(n6160), .ZN(n2460) );
  NAND2_X1 U1215 ( .A1(n2333), .A2(n3892), .ZN(n297) );
  NAND2_X2 U1217 ( .A1(n298), .A2(n297), .ZN(n3856) );
  INV_X1 U1219 ( .A(n3892), .ZN(n296) );
  NAND2_X2 U1222 ( .A1(n300), .A2(n301), .ZN(n303) );
  OAI21_X2 U1225 ( .B1(n3075), .B2(n3076), .A(n6587), .ZN(n1181) );
  MUX2_X2 U1229 ( .A(n6029), .B(n5895), .S(b[0]), .Z(n4437) );
  NAND2_X1 U1232 ( .A1(n3942), .A2(n2587), .ZN(n307) );
  NAND2_X2 U1233 ( .A1(n305), .A2(n306), .ZN(n308) );
  NAND2_X2 U1234 ( .A1(n307), .A2(n308), .ZN(n3976) );
  INV_X2 U1235 ( .A(n3942), .ZN(n305) );
  INV_X2 U1236 ( .A(n2587), .ZN(n306) );
  INV_X1 U1239 ( .A(n4939), .ZN(n1479) );
  XNOR2_X2 U1240 ( .A(n4315), .B(n4314), .ZN(n1431) );
  INV_X8 U1245 ( .A(a[16]), .ZN(n311) );
  XOR2_X2 U1247 ( .A(a[3]), .B(b[20]), .Z(n2743) );
  NAND2_X1 U1250 ( .A1(n1565), .A2(n4447), .ZN(n317) );
  NAND2_X2 U1252 ( .A1(n317), .A2(n318), .ZN(n4466) );
  INV_X8 U1257 ( .A(b[23]), .ZN(n1075) );
  OAI22_X1 U1258 ( .A1(n3959), .A2(n4689), .B1(n3958), .B2(b[9]), .ZN(n3961)
         );
  NAND2_X1 U1259 ( .A1(n4689), .A2(b[19]), .ZN(n3683) );
  NAND2_X1 U1261 ( .A1(n432), .A2(n2929), .ZN(n319) );
  NAND2_X4 U1262 ( .A1(n4899), .A2(n689), .ZN(n432) );
  NAND2_X2 U1265 ( .A1(n2987), .A2(n2373), .ZN(n320) );
  NAND2_X2 U1266 ( .A1(n3008), .A2(n4009), .ZN(n538) );
  NAND2_X1 U1269 ( .A1(n4998), .A2(n4392), .ZN(n4394) );
  NAND2_X2 U1270 ( .A1(n3308), .A2(n2738), .ZN(n3700) );
  XOR2_X2 U1271 ( .A(n4056), .B(n4061), .Z(n3945) );
  NOR2_X2 U1272 ( .A1(n3938), .A2(n3654), .ZN(n1914) );
  INV_X4 U1273 ( .A(n2300), .ZN(n809) );
  INV_X4 U1274 ( .A(n2031), .ZN(n321) );
  AOI22_X2 U1276 ( .A1(n2803), .A2(n1006), .B1(n2803), .B2(n3408), .ZN(n324)
         );
  NOR2_X4 U1277 ( .A1(n3235), .A2(n3234), .ZN(n3408) );
  OAI21_X2 U1278 ( .B1(n4484), .B2(n3051), .A(n1004), .ZN(n2403) );
  NAND2_X2 U1280 ( .A1(n1826), .A2(n1825), .ZN(n326) );
  INV_X1 U1283 ( .A(n2391), .ZN(n1082) );
  NAND2_X1 U1284 ( .A1(n4219), .A2(n2249), .ZN(n4131) );
  AOI22_X1 U1286 ( .A1(a[0]), .A2(n4188), .B1(n4219), .B2(n3342), .ZN(n4189)
         );
  NAND2_X4 U1289 ( .A1(n5070), .A2(a[19]), .ZN(n328) );
  NAND2_X1 U1290 ( .A1(n5287), .A2(n5355), .ZN(n331) );
  NAND2_X2 U1291 ( .A1(n329), .A2(n330), .ZN(n332) );
  NAND2_X2 U1292 ( .A1(n331), .A2(n332), .ZN(n5331) );
  INV_X2 U1293 ( .A(n5287), .ZN(n329) );
  INV_X1 U1294 ( .A(n5355), .ZN(n330) );
  NOR2_X2 U1296 ( .A1(n3704), .A2(n4704), .ZN(n1790) );
  NAND2_X1 U1297 ( .A1(b[21]), .A2(n3581), .ZN(n3600) );
  NOR2_X2 U1298 ( .A1(n4919), .A2(n3575), .ZN(n2752) );
  NOR2_X4 U1299 ( .A1(n4979), .A2(n4976), .ZN(n5851) );
  AOI22_X2 U1300 ( .A1(n4780), .A2(n3313), .B1(n1440), .B2(n4779), .ZN(n4962)
         );
  INV_X1 U1301 ( .A(n3900), .ZN(n3886) );
  NOR2_X1 U1304 ( .A1(n5149), .A2(n2358), .ZN(n2357) );
  OAI21_X1 U1305 ( .B1(n2489), .B2(n5149), .A(n2358), .ZN(n2355) );
  NAND2_X2 U1306 ( .A1(n333), .A2(n334), .ZN(n336) );
  INV_X4 U1310 ( .A(n4034), .ZN(n4038) );
  NAND2_X1 U1312 ( .A1(n4504), .A2(b[18]), .ZN(n3329) );
  NOR2_X2 U1315 ( .A1(n4499), .A2(n4498), .ZN(n3430) );
  NAND2_X4 U1318 ( .A1(n338), .A2(n339), .ZN(n3190) );
  INV_X8 U1320 ( .A(b[5]), .ZN(n3870) );
  NOR2_X1 U1321 ( .A1(n1012), .A2(b[12]), .ZN(n1735) );
  NAND2_X2 U1322 ( .A1(n4933), .A2(n4811), .ZN(n1504) );
  NAND2_X2 U1324 ( .A1(n1019), .A2(n5307), .ZN(n5317) );
  NAND2_X2 U1325 ( .A1(n1240), .A2(n4901), .ZN(n340) );
  NAND2_X2 U1326 ( .A1(n2251), .A2(n2254), .ZN(n341) );
  NAND2_X1 U1329 ( .A1(n4370), .A2(n3695), .ZN(n342) );
  NAND2_X2 U1330 ( .A1(n881), .A2(n4976), .ZN(n343) );
  NOR3_X4 U1334 ( .A1(n1609), .A2(n1610), .A3(n5572), .ZN(n5913) );
  NAND2_X2 U1335 ( .A1(n1099), .A2(n5384), .ZN(n345) );
  NAND2_X1 U1338 ( .A1(n1776), .A2(n4457), .ZN(n349) );
  INV_X2 U1339 ( .A(n1776), .ZN(n347) );
  INV_X1 U1345 ( .A(n4019), .ZN(n351) );
  OAI21_X1 U1346 ( .B1(n4289), .B2(n4288), .A(n4287), .ZN(n4302) );
  INV_X2 U1350 ( .A(n4903), .ZN(n354) );
  NAND2_X4 U1351 ( .A1(a[10]), .A2(a[9]), .ZN(n360) );
  NAND2_X2 U1352 ( .A1(n466), .A2(n359), .ZN(n361) );
  INV_X8 U1355 ( .A(a[9]), .ZN(n359) );
  OAI21_X2 U1359 ( .B1(n1721), .B2(n1720), .A(n5564), .ZN(n1719) );
  NAND2_X4 U1360 ( .A1(a[2]), .A2(a[1]), .ZN(n365) );
  NAND2_X2 U1361 ( .A1(n672), .A2(n673), .ZN(n366) );
  NOR2_X1 U1362 ( .A1(n1000), .A2(n367), .ZN(n947) );
  NAND2_X1 U1363 ( .A1(a[11]), .A2(n3154), .ZN(n367) );
  NAND2_X2 U1364 ( .A1(n1261), .A2(n1260), .ZN(n368) );
  NAND2_X2 U1365 ( .A1(n5610), .A2(n5609), .ZN(n5888) );
  NAND2_X1 U1366 ( .A1(n1716), .A2(n1715), .ZN(n372) );
  NAND2_X2 U1367 ( .A1(n370), .A2(n371), .ZN(n373) );
  NAND2_X2 U1368 ( .A1(n373), .A2(n372), .ZN(n1714) );
  INV_X2 U1369 ( .A(n1716), .ZN(n370) );
  INV_X2 U1370 ( .A(n1715), .ZN(n371) );
  NAND2_X1 U1371 ( .A1(n2629), .A2(n2066), .ZN(n376) );
  NAND2_X2 U1372 ( .A1(n374), .A2(n375), .ZN(n377) );
  NAND2_X2 U1373 ( .A1(n376), .A2(n377), .ZN(n4871) );
  INV_X4 U1374 ( .A(n2629), .ZN(n374) );
  INV_X2 U1375 ( .A(n2066), .ZN(n375) );
  NAND2_X1 U1378 ( .A1(n2651), .A2(n4452), .ZN(n380) );
  INV_X2 U1381 ( .A(n2651), .ZN(n378) );
  AOI21_X2 U1383 ( .B1(n2326), .B2(n4025), .A(n1874), .ZN(n4452) );
  NAND3_X2 U1384 ( .A1(n3338), .A2(n3337), .A3(n4628), .ZN(n3336) );
  NAND2_X1 U1385 ( .A1(n2537), .A2(b[19]), .ZN(n383) );
  NAND2_X1 U1386 ( .A1(n3438), .A2(n5266), .ZN(n384) );
  NAND2_X1 U1389 ( .A1(n5459), .A2(n5458), .ZN(n386) );
  NAND2_X2 U1390 ( .A1(n385), .A2(n1344), .ZN(n387) );
  NOR2_X2 U1392 ( .A1(n2331), .A2(n2330), .ZN(n2329) );
  NAND2_X1 U1393 ( .A1(n5298), .A2(n5303), .ZN(n391) );
  NAND2_X1 U1396 ( .A1(n1406), .A2(n5297), .ZN(n394) );
  NAND2_X4 U1399 ( .A1(a[22]), .A2(a[21]), .ZN(n395) );
  XNOR2_X2 U1404 ( .A(b[6]), .B(a[21]), .ZN(n4703) );
  XNOR2_X2 U1405 ( .A(b[12]), .B(a[21]), .ZN(n4994) );
  XNOR2_X2 U1406 ( .A(a[21]), .B(b[1]), .ZN(n4434) );
  INV_X8 U1407 ( .A(a[21]), .ZN(n4989) );
  INV_X1 U1409 ( .A(n2809), .ZN(n489) );
  NOR2_X2 U1410 ( .A1(n3916), .A2(n3917), .ZN(n2809) );
  INV_X1 U1415 ( .A(n4568), .ZN(n4569) );
  INV_X4 U1416 ( .A(n5084), .ZN(n1830) );
  INV_X1 U1417 ( .A(n2594), .ZN(n1800) );
  OAI21_X1 U1419 ( .B1(n5024), .B2(n985), .A(n3088), .ZN(n2397) );
  NAND2_X2 U1421 ( .A1(n5176), .A2(n2401), .ZN(n1629) );
  INV_X4 U1424 ( .A(n1765), .ZN(n397) );
  INV_X1 U1426 ( .A(n3981), .ZN(n3982) );
  INV_X1 U1427 ( .A(n3923), .ZN(n2843) );
  NOR2_X1 U1429 ( .A1(n3323), .A2(n4769), .ZN(n400) );
  NOR2_X2 U1430 ( .A1(n3323), .A2(n4769), .ZN(n401) );
  NOR2_X4 U1432 ( .A1(n4407), .A2(n4406), .ZN(n4413) );
  NAND2_X1 U1434 ( .A1(n3919), .A2(n4059), .ZN(n405) );
  NAND2_X2 U1435 ( .A1(n3943), .A2(n4065), .ZN(n406) );
  NAND2_X2 U1436 ( .A1(n405), .A2(n406), .ZN(n3166) );
  NAND2_X2 U1439 ( .A1(n2010), .A2(n2322), .ZN(n3939) );
  INV_X1 U1440 ( .A(n3943), .ZN(n3919) );
  NAND2_X1 U1442 ( .A1(n1746), .A2(n5155), .ZN(n409) );
  NAND2_X2 U1443 ( .A1(n407), .A2(n408), .ZN(n410) );
  NAND2_X2 U1444 ( .A1(n409), .A2(n410), .ZN(n3403) );
  INV_X2 U1445 ( .A(n1746), .ZN(n407) );
  INV_X1 U1446 ( .A(n5155), .ZN(n408) );
  NAND2_X1 U1447 ( .A1(n2537), .A2(b[14]), .ZN(n412) );
  NAND2_X1 U1448 ( .A1(n5293), .A2(n5266), .ZN(n413) );
  NAND2_X2 U1449 ( .A1(n412), .A2(n413), .ZN(n5072) );
  INV_X4 U1451 ( .A(n4408), .ZN(n414) );
  INV_X4 U1452 ( .A(n4408), .ZN(n1455) );
  NOR2_X1 U1453 ( .A1(n4058), .A2(n4064), .ZN(n3944) );
  NAND2_X4 U1455 ( .A1(n1259), .A2(n1258), .ZN(n1148) );
  NAND2_X2 U1456 ( .A1(n6214), .A2(n1041), .ZN(n415) );
  INV_X4 U1458 ( .A(n1484), .ZN(n4524) );
  INV_X4 U1459 ( .A(n5457), .ZN(n416) );
  NAND2_X2 U1461 ( .A1(n2102), .A2(n3492), .ZN(n2690) );
  INV_X1 U1465 ( .A(n4914), .ZN(n418) );
  NAND2_X2 U1466 ( .A1(n3468), .A2(n2613), .ZN(n584) );
  NOR2_X1 U1467 ( .A1(n5672), .A2(n3722), .ZN(n421) );
  BUF_X4 U1468 ( .A(n5667), .Z(n422) );
  NOR2_X2 U1469 ( .A1(n4099), .A2(n424), .ZN(n425) );
  INV_X4 U1472 ( .A(n4100), .ZN(n424) );
  NAND2_X1 U1477 ( .A1(n3409), .A2(n2929), .ZN(n434) );
  NOR2_X4 U1478 ( .A1(n4845), .A2(n5952), .ZN(n430) );
  AOI21_X1 U1480 ( .B1(b[5]), .B2(n4812), .A(a[23]), .ZN(n4814) );
  NAND2_X2 U1481 ( .A1(n581), .A2(n830), .ZN(n832) );
  NAND2_X2 U1482 ( .A1(n4856), .A2(n4863), .ZN(n1556) );
  NOR2_X2 U1483 ( .A1(n3461), .A2(n5707), .ZN(n3362) );
  NOR2_X2 U1485 ( .A1(n2249), .A2(n1194), .ZN(n4050) );
  INV_X4 U1486 ( .A(n4442), .ZN(n3331) );
  NAND3_X1 U1488 ( .A1(n6015), .A2(n6014), .A3(n3476), .ZN(n6019) );
  NAND2_X1 U1491 ( .A1(n2230), .A2(n2231), .ZN(n1545) );
  NAND2_X1 U1492 ( .A1(n4219), .A2(n4942), .ZN(n3994) );
  NOR2_X1 U1493 ( .A1(n5620), .A2(n5377), .ZN(n6016) );
  NAND2_X1 U1494 ( .A1(n2724), .A2(n4408), .ZN(n470) );
  NAND2_X1 U1495 ( .A1(n4775), .A2(n6654), .ZN(n3204) );
  NAND2_X2 U1496 ( .A1(a[23]), .A2(n2038), .ZN(n435) );
  INV_X1 U1499 ( .A(n4921), .ZN(n493) );
  NAND2_X1 U1501 ( .A1(n868), .A2(n869), .ZN(n716) );
  NAND2_X1 U1503 ( .A1(n434), .A2(n432), .ZN(n437) );
  INV_X1 U1504 ( .A(n2235), .ZN(n438) );
  NOR2_X2 U1507 ( .A1(a[11]), .A2(n468), .ZN(n441) );
  INV_X4 U1508 ( .A(n4295), .ZN(n3289) );
  NOR2_X4 U1509 ( .A1(n817), .A2(n3540), .ZN(n3831) );
  INV_X1 U1512 ( .A(n3283), .ZN(n650) );
  NAND3_X2 U1513 ( .A1(n4966), .A2(n5092), .A3(n2928), .ZN(n3370) );
  NAND2_X2 U1514 ( .A1(n2853), .A2(n6596), .ZN(n1071) );
  NOR2_X1 U1516 ( .A1(n1023), .A2(n5332), .ZN(n5334) );
  INV_X4 U1518 ( .A(n2099), .ZN(n446) );
  NOR3_X1 U1519 ( .A1(n1996), .A2(n4650), .A3(n4651), .ZN(n1991) );
  NAND2_X2 U1521 ( .A1(n1596), .A2(n1595), .ZN(n452) );
  INV_X1 U1522 ( .A(n3108), .ZN(n1379) );
  NOR2_X4 U1523 ( .A1(n3817), .A2(n3816), .ZN(n3820) );
  NOR2_X2 U1524 ( .A1(n3815), .A2(n3617), .ZN(n3817) );
  NAND2_X4 U1531 ( .A1(n2151), .A2(n2153), .ZN(n4974) );
  NAND2_X2 U1532 ( .A1(n821), .A2(n822), .ZN(n824) );
  NOR2_X4 U1533 ( .A1(n327), .A2(n4413), .ZN(n458) );
  INV_X4 U1534 ( .A(n458), .ZN(n3570) );
  AOI21_X1 U1535 ( .B1(n5876), .B2(n5862), .A(n5875), .ZN(n5868) );
  BUF_X4 U1537 ( .A(n4874), .Z(n459) );
  INV_X1 U1538 ( .A(n4630), .ZN(n3337) );
  NAND2_X2 U1539 ( .A1(n4863), .A2(n4866), .ZN(n2639) );
  INV_X4 U1540 ( .A(n460), .ZN(n3867) );
  NAND2_X4 U1542 ( .A1(n1436), .A2(n4657), .ZN(n1387) );
  INV_X8 U1546 ( .A(a[8]), .ZN(n4389) );
  NAND2_X2 U1547 ( .A1(a[9]), .A2(n4389), .ZN(n3958) );
  INV_X4 U1548 ( .A(n461), .ZN(n531) );
  NOR2_X2 U1549 ( .A1(n4995), .A2(b[8]), .ZN(n463) );
  INV_X4 U1551 ( .A(n5840), .ZN(n1274) );
  NAND2_X2 U1553 ( .A1(n1510), .A2(n1509), .ZN(n753) );
  INV_X1 U1554 ( .A(n5610), .ZN(n5611) );
  NOR2_X2 U1555 ( .A1(n5453), .A2(n5452), .ZN(n5553) );
  INV_X4 U1558 ( .A(n5999), .ZN(n1607) );
  NOR2_X1 U1559 ( .A1(n5491), .A2(n5490), .ZN(n5493) );
  NAND2_X2 U1560 ( .A1(n754), .A2(n755), .ZN(n757) );
  NAND2_X4 U1562 ( .A1(a[10]), .A2(a[9]), .ZN(n468) );
  NOR2_X2 U1567 ( .A1(n2889), .A2(n4342), .ZN(n3050) );
  NAND2_X2 U1568 ( .A1(n2724), .A2(n4408), .ZN(n3736) );
  NAND2_X1 U1570 ( .A1(a[1]), .A2(n2563), .ZN(n471) );
  NAND2_X1 U1571 ( .A1(a[1]), .A2(n2563), .ZN(n472) );
  NOR2_X4 U1574 ( .A1(n2054), .A2(n2811), .ZN(n5368) );
  NOR2_X4 U1576 ( .A1(n6504), .A2(n3355), .ZN(n4309) );
  INV_X4 U1577 ( .A(n2927), .ZN(n2918) );
  INV_X8 U1578 ( .A(a[12]), .ZN(n3792) );
  INV_X4 U1580 ( .A(n4601), .ZN(n4506) );
  NOR2_X4 U1581 ( .A1(n2199), .A2(n2198), .ZN(n3887) );
  AOI22_X2 U1582 ( .A1(n4774), .A2(b[2]), .B1(n2249), .B2(n699), .ZN(n2198) );
  OAI21_X2 U1583 ( .B1(n3935), .B2(n3936), .A(n3934), .ZN(n3983) );
  NAND2_X2 U1584 ( .A1(n588), .A2(n4654), .ZN(n591) );
  INV_X1 U1585 ( .A(n4917), .ZN(n2758) );
  NAND2_X2 U1588 ( .A1(n2516), .A2(n283), .ZN(n2515) );
  NOR2_X4 U1590 ( .A1(n2830), .A2(n2603), .ZN(n2310) );
  NAND2_X2 U1591 ( .A1(n1544), .A2(n1543), .ZN(n477) );
  NAND2_X2 U1594 ( .A1(n3695), .A2(n4370), .ZN(n4372) );
  NAND2_X1 U1595 ( .A1(n3088), .A2(n985), .ZN(n480) );
  NAND2_X2 U1596 ( .A1(n478), .A2(n479), .ZN(n481) );
  NAND2_X2 U1597 ( .A1(n480), .A2(n481), .ZN(n2300) );
  AOI21_X2 U1600 ( .B1(n5451), .B2(n5450), .A(n5449), .ZN(n5453) );
  NAND2_X2 U1602 ( .A1(n2600), .A2(n2599), .ZN(n482) );
  NAND2_X2 U1603 ( .A1(n2303), .A2(n557), .ZN(n483) );
  NAND2_X2 U1604 ( .A1(n557), .A2(n2303), .ZN(n484) );
  OAI22_X1 U1607 ( .A1(n6031), .A2(n6030), .B1(n6029), .B2(n6028), .ZN(n6122)
         );
  INV_X1 U1608 ( .A(n4479), .ZN(n4473) );
  NAND2_X2 U1611 ( .A1(n5035), .A2(n556), .ZN(n5036) );
  NOR2_X4 U1613 ( .A1(n2918), .A2(n2917), .ZN(n2925) );
  NAND3_X2 U1614 ( .A1(n4490), .A2(n5529), .A3(a[1]), .ZN(n2923) );
  INV_X1 U1616 ( .A(n5888), .ZN(n5916) );
  NAND2_X4 U1617 ( .A1(n5678), .A2(n3453), .ZN(n3153) );
  INV_X1 U1618 ( .A(n4901), .ZN(n3188) );
  NAND2_X1 U1619 ( .A1(n647), .A2(n1263), .ZN(n486) );
  NAND2_X1 U1620 ( .A1(n441), .A2(b[4]), .ZN(n2196) );
  NAND2_X1 U1623 ( .A1(n3166), .A2(n2809), .ZN(n490) );
  NAND2_X2 U1624 ( .A1(n488), .A2(n489), .ZN(n491) );
  INV_X2 U1626 ( .A(n3166), .ZN(n488) );
  INV_X4 U1627 ( .A(n3011), .ZN(n3586) );
  NAND2_X2 U1629 ( .A1(n747), .A2(n761), .ZN(n750) );
  INV_X1 U1630 ( .A(n3545), .ZN(n522) );
  NAND2_X1 U1631 ( .A1(n4920), .A2(n4921), .ZN(n494) );
  INV_X1 U1633 ( .A(n4920), .ZN(n492) );
  NAND2_X2 U1636 ( .A1(n5059), .A2(n5117), .ZN(n831) );
  BUF_X4 U1637 ( .A(n5566), .Z(n3160) );
  NAND2_X1 U1640 ( .A1(n5451), .A2(n2870), .ZN(n499) );
  INV_X2 U1644 ( .A(n2870), .ZN(n498) );
  NAND2_X2 U1647 ( .A1(n503), .A2(n504), .ZN(n1978) );
  INV_X8 U1648 ( .A(a[14]), .ZN(n501) );
  INV_X8 U1649 ( .A(a[13]), .ZN(n502) );
  INV_X1 U1650 ( .A(n4078), .ZN(n4080) );
  NAND3_X2 U1651 ( .A1(n4863), .A2(n4865), .A3(n4864), .ZN(n2640) );
  NOR2_X4 U1653 ( .A1(a[4]), .A2(a[3]), .ZN(n505) );
  NOR2_X4 U1654 ( .A1(a[4]), .A2(a[3]), .ZN(n506) );
  NAND2_X2 U1655 ( .A1(n2152), .A2(n6093), .ZN(n2151) );
  INV_X4 U1656 ( .A(n3190), .ZN(n2110) );
  NAND2_X2 U1657 ( .A1(n507), .A2(n508), .ZN(n510) );
  NAND2_X1 U1659 ( .A1(n816), .A2(n815), .ZN(n511) );
  OAI21_X2 U1661 ( .B1(n5079), .B2(n5220), .A(n3504), .ZN(n5295) );
  NOR3_X4 U1663 ( .A1(n3684), .A2(a[7]), .A3(a[8]), .ZN(n512) );
  NOR3_X4 U1664 ( .A1(n3684), .A2(a[7]), .A3(a[8]), .ZN(n513) );
  NAND2_X2 U1668 ( .A1(n515), .A2(n514), .ZN(n517) );
  NAND2_X2 U1673 ( .A1(n518), .A2(n519), .ZN(n521) );
  INV_X1 U1674 ( .A(n4867), .ZN(n519) );
  NAND2_X1 U1675 ( .A1(n523), .A2(n3545), .ZN(n524) );
  NAND2_X2 U1676 ( .A1(n522), .A2(n4763), .ZN(n525) );
  INV_X2 U1677 ( .A(n4763), .ZN(n523) );
  XOR2_X2 U1681 ( .A(b[9]), .B(a[19]), .Z(n530) );
  NAND2_X1 U1686 ( .A1(n2267), .A2(n2268), .ZN(n710) );
  NOR2_X1 U1689 ( .A1(n2155), .A2(n2086), .ZN(n5828) );
  NAND2_X1 U1690 ( .A1(n2200), .A2(n2201), .ZN(n1299) );
  NAND2_X1 U1691 ( .A1(n4598), .A2(n267), .ZN(n1886) );
  NOR2_X1 U1692 ( .A1(n1847), .A2(b[1]), .ZN(n1768) );
  NAND2_X1 U1693 ( .A1(n4475), .A2(n4474), .ZN(n536) );
  NAND2_X2 U1695 ( .A1(n537), .A2(n536), .ZN(n1110) );
  NAND2_X2 U1697 ( .A1(n2638), .A2(n6325), .ZN(n2637) );
  NAND2_X1 U1699 ( .A1(n1435), .A2(n3894), .ZN(n1434) );
  NAND2_X2 U1700 ( .A1(n5342), .A2(n5341), .ZN(n5451) );
  NOR2_X2 U1701 ( .A1(n1153), .A2(n1154), .ZN(n539) );
  NOR2_X2 U1702 ( .A1(n1154), .A2(n1153), .ZN(n2865) );
  NAND2_X1 U1704 ( .A1(b[12]), .A2(n4601), .ZN(n1927) );
  OR2_X4 U1705 ( .A1(n3465), .A2(n4601), .ZN(n2746) );
  NAND2_X1 U1706 ( .A1(b[16]), .A2(n4601), .ZN(n2161) );
  NOR2_X1 U1707 ( .A1(n3540), .A2(n4601), .ZN(n1920) );
  NAND2_X4 U1708 ( .A1(n3239), .A2(n3063), .ZN(n4581) );
  AOI21_X1 U1710 ( .B1(n5376), .B2(n5621), .A(n5620), .ZN(n5390) );
  INV_X1 U1711 ( .A(n1840), .ZN(n5792) );
  NAND2_X2 U1712 ( .A1(n5074), .A2(n3367), .ZN(n1687) );
  NAND2_X1 U1714 ( .A1(n4194), .A2(n2339), .ZN(n542) );
  INV_X2 U1717 ( .A(n4194), .ZN(n540) );
  INV_X2 U1718 ( .A(n2339), .ZN(n541) );
  NAND2_X1 U1719 ( .A1(n1633), .A2(n4205), .ZN(n546) );
  INV_X2 U1722 ( .A(n1633), .ZN(n544) );
  NAND2_X1 U1724 ( .A1(n1137), .A2(n1136), .ZN(n549) );
  NAND2_X2 U1725 ( .A1(n549), .A2(n550), .ZN(n5676) );
  INV_X2 U1726 ( .A(n1137), .ZN(n548) );
  NAND2_X1 U1727 ( .A1(n2519), .A2(n102), .ZN(n553) );
  NAND2_X2 U1728 ( .A1(n551), .A2(n552), .ZN(n554) );
  NAND2_X2 U1729 ( .A1(n553), .A2(n554), .ZN(n1137) );
  INV_X2 U1730 ( .A(n2519), .ZN(n551) );
  INV_X1 U1733 ( .A(n5031), .ZN(n556) );
  NAND3_X2 U1736 ( .A1(n563), .A2(n6607), .A3(n4642), .ZN(n2039) );
  INV_X4 U1739 ( .A(n5040), .ZN(n1941) );
  INV_X1 U1740 ( .A(n3431), .ZN(n975) );
  NAND2_X2 U1741 ( .A1(n559), .A2(n560), .ZN(n562) );
  AOI22_X1 U1746 ( .A1(n4662), .A2(n2967), .B1(n4661), .B2(n2695), .ZN(n4720)
         );
  NAND2_X2 U1747 ( .A1(n1059), .A2(n4586), .ZN(n2967) );
  NAND2_X1 U1750 ( .A1(n1083), .A2(n1628), .ZN(n571) );
  NAND2_X2 U1752 ( .A1(n571), .A2(n572), .ZN(n2391) );
  NAND2_X1 U1754 ( .A1(n4917), .A2(n4916), .ZN(n575) );
  NAND2_X2 U1755 ( .A1(n573), .A2(n574), .ZN(n576) );
  NOR2_X1 U1757 ( .A1(n2327), .A2(n4997), .ZN(n3631) );
  XNOR2_X2 U1764 ( .A(n2512), .B(n4046), .ZN(n581) );
  INV_X4 U1765 ( .A(n581), .ZN(n5059) );
  NAND2_X2 U1766 ( .A1(n3620), .A2(n3083), .ZN(n2902) );
  OAI22_X2 U1767 ( .A1(n2129), .A2(b[18]), .B1(n648), .B2(n5529), .ZN(n2128)
         );
  NAND2_X4 U1768 ( .A1(n1360), .A2(n2124), .ZN(n2131) );
  NAND2_X1 U1772 ( .A1(n1549), .A2(n3996), .ZN(n1553) );
  NAND2_X1 U1773 ( .A1(n1550), .A2(n3996), .ZN(n1871) );
  AOI22_X2 U1774 ( .A1(n6569), .A2(n4795), .B1(n606), .B2(b[1]), .ZN(n4211) );
  INV_X4 U1775 ( .A(n3492), .ZN(n2101) );
  NAND2_X2 U1776 ( .A1(n2435), .A2(n2434), .ZN(n585) );
  NAND2_X2 U1777 ( .A1(n2435), .A2(n2434), .ZN(n586) );
  NAND2_X4 U1781 ( .A1(n2699), .A2(a[19]), .ZN(n2434) );
  NAND2_X2 U1783 ( .A1(n2818), .A2(n4668), .ZN(n2968) );
  NAND2_X2 U1785 ( .A1(n6204), .A2(n593), .ZN(n595) );
  INV_X2 U1787 ( .A(n3313), .ZN(n593) );
  NAND2_X1 U1788 ( .A1(n401), .A2(n4802), .ZN(n598) );
  NAND2_X2 U1790 ( .A1(n598), .A2(n599), .ZN(n3150) );
  INV_X4 U1794 ( .A(n2336), .ZN(n4606) );
  NAND2_X2 U1795 ( .A1(n5384), .A2(n1099), .ZN(n600) );
  NAND2_X2 U1796 ( .A1(n646), .A2(n3500), .ZN(n601) );
  NAND2_X1 U1801 ( .A1(n2082), .A2(n2676), .ZN(n604) );
  NAND2_X2 U1802 ( .A1(n602), .A2(n603), .ZN(n605) );
  INV_X2 U1803 ( .A(n2082), .ZN(n602) );
  INV_X1 U1804 ( .A(n2676), .ZN(n603) );
  NAND2_X2 U1805 ( .A1(n6207), .A2(n1870), .ZN(n3315) );
  INV_X1 U1806 ( .A(n5817), .ZN(n2154) );
  NAND2_X1 U1807 ( .A1(n998), .A2(n6221), .ZN(n1104) );
  NAND2_X2 U1808 ( .A1(n2300), .A2(n5023), .ZN(n811) );
  NOR2_X2 U1809 ( .A1(n5888), .A2(n5875), .ZN(n6005) );
  NOR2_X4 U1810 ( .A1(n3305), .A2(a[9]), .ZN(n606) );
  NAND2_X2 U1812 ( .A1(n4746), .A2(n5277), .ZN(n4348) );
  INV_X4 U1814 ( .A(n4549), .ZN(n608) );
  NAND2_X2 U1815 ( .A1(n4554), .A2(n4555), .ZN(n2806) );
  NAND2_X2 U1816 ( .A1(n1882), .A2(n1881), .ZN(n4554) );
  AND2_X2 U1817 ( .A1(n609), .A2(n585), .ZN(n2253) );
  XOR2_X2 U1818 ( .A(b[9]), .B(a[21]), .Z(n609) );
  INV_X4 U1819 ( .A(n5072), .ZN(n3450) );
  NOR2_X2 U1820 ( .A1(n3622), .A2(n5072), .ZN(n2354) );
  OAI21_X2 U1821 ( .B1(n1875), .B2(n1813), .A(n1805), .ZN(n1812) );
  NAND2_X1 U1822 ( .A1(n4566), .A2(n4568), .ZN(n4570) );
  NAND2_X2 U1826 ( .A1(n1149), .A2(n4232), .ZN(n1152) );
  NAND2_X2 U1828 ( .A1(n2510), .A2(n4942), .ZN(n3296) );
  INV_X4 U1829 ( .A(n5374), .ZN(n3663) );
  INV_X1 U1830 ( .A(n5853), .ZN(n3389) );
  INV_X4 U1834 ( .A(n1148), .ZN(n4763) );
  XOR2_X2 U1835 ( .A(a[21]), .B(b[3]), .Z(n611) );
  INV_X8 U1837 ( .A(n4483), .ZN(n2950) );
  INV_X4 U1844 ( .A(n4232), .ZN(n1151) );
  OAI21_X1 U1845 ( .B1(n5660), .B2(n4150), .A(n4149), .ZN(n688) );
  NAND2_X4 U1849 ( .A1(n1978), .A2(a[15]), .ZN(n2932) );
  NAND2_X2 U1851 ( .A1(n614), .A2(n615), .ZN(n3746) );
  NOR2_X2 U1855 ( .A1(n6331), .A2(n5383), .ZN(n616) );
  NOR2_X1 U1856 ( .A1(n2517), .A2(n1031), .ZN(n1505) );
  NAND2_X1 U1857 ( .A1(n1120), .A2(n2438), .ZN(n619) );
  NAND2_X2 U1858 ( .A1(n617), .A2(n618), .ZN(n620) );
  INV_X2 U1859 ( .A(n1120), .ZN(n617) );
  INV_X2 U1860 ( .A(n2438), .ZN(n618) );
  NOR2_X2 U1861 ( .A1(n5276), .A2(n5275), .ZN(n5345) );
  NAND2_X1 U1865 ( .A1(n465), .A2(b[13]), .ZN(n3691) );
  OAI21_X2 U1866 ( .B1(n4633), .B2(n4632), .A(n4631), .ZN(n1076) );
  AOI21_X1 U1867 ( .B1(n4404), .B2(n6610), .A(n4402), .ZN(n4523) );
  NOR2_X2 U1869 ( .A1(n3622), .A2(n5072), .ZN(n5112) );
  NOR2_X4 U1871 ( .A1(n999), .A2(a[11]), .ZN(n3581) );
  NAND2_X1 U1876 ( .A1(n1622), .A2(n1674), .ZN(n626) );
  NAND2_X4 U1878 ( .A1(n626), .A2(n627), .ZN(n5472) );
  INV_X2 U1879 ( .A(n1622), .ZN(n624) );
  INV_X4 U1880 ( .A(n1674), .ZN(n625) );
  INV_X4 U1882 ( .A(n5472), .ZN(n5525) );
  INV_X4 U1883 ( .A(n3620), .ZN(n1709) );
  NOR2_X4 U1884 ( .A1(n5377), .A2(n616), .ZN(n628) );
  OAI21_X2 U1885 ( .B1(n951), .B2(n436), .A(n1660), .ZN(n629) );
  OAI21_X1 U1886 ( .B1(n951), .B2(n436), .A(n1660), .ZN(n4959) );
  NAND2_X2 U1888 ( .A1(n749), .A2(n750), .ZN(n5172) );
  OAI22_X2 U1889 ( .A1(n5991), .A2(n1013), .B1(n5983), .B2(n5982), .ZN(n5989)
         );
  INV_X1 U1890 ( .A(n4373), .ZN(n3738) );
  BUF_X4 U1891 ( .A(n4969), .Z(n630) );
  NAND2_X2 U1893 ( .A1(n1844), .A2(n2488), .ZN(n2837) );
  NAND2_X1 U1894 ( .A1(b[6]), .A2(n5218), .ZN(n4320) );
  NAND2_X2 U1898 ( .A1(n4731), .A2(n4730), .ZN(n1483) );
  NOR2_X2 U1899 ( .A1(n2587), .A2(n3942), .ZN(n4061) );
  NAND2_X2 U1901 ( .A1(n934), .A2(n933), .ZN(n4838) );
  OAI21_X1 U1905 ( .B1(n5217), .B2(n5206), .A(n5216), .ZN(n637) );
  OAI21_X1 U1908 ( .B1(n5206), .B2(n5217), .A(n5216), .ZN(n5630) );
  OAI22_X2 U1909 ( .A1(n5120), .A2(n2512), .B1(n5119), .B2(n5118), .ZN(n5177)
         );
  NAND2_X1 U1910 ( .A1(n2538), .A2(n2539), .ZN(n642) );
  NAND2_X2 U1911 ( .A1(n640), .A2(n641), .ZN(n643) );
  NAND2_X2 U1912 ( .A1(n643), .A2(n642), .ZN(n5780) );
  NAND2_X4 U1915 ( .A1(n4601), .A2(b[14]), .ZN(n646) );
  NOR2_X1 U1917 ( .A1(n3831), .A2(n3833), .ZN(n3029) );
  INV_X4 U1919 ( .A(n5077), .ZN(n5336) );
  NOR2_X4 U1922 ( .A1(n1745), .A2(n1744), .ZN(n5383) );
  OAI21_X1 U1924 ( .B1(n2195), .B2(n3887), .A(n2437), .ZN(n766) );
  INV_X4 U1927 ( .A(n4070), .ZN(n4072) );
  NOR2_X4 U1928 ( .A1(n3913), .A2(n2974), .ZN(n4070) );
  NOR2_X2 U1931 ( .A1(n5105), .A2(n6527), .ZN(n1988) );
  NAND3_X1 U1932 ( .A1(n943), .A2(n4511), .A3(n4510), .ZN(n2788) );
  NAND2_X2 U1933 ( .A1(n3201), .A2(n2913), .ZN(n647) );
  AOI22_X2 U1935 ( .A1(b[19]), .A2(n4405), .B1(n3438), .B2(n1012), .ZN(n4407)
         );
  NAND2_X4 U1936 ( .A1(n1946), .A2(n995), .ZN(n3318) );
  INV_X4 U1939 ( .A(n5897), .ZN(n3351) );
  NAND3_X1 U1940 ( .A1(n4219), .A2(n3465), .A3(n3540), .ZN(n2096) );
  XNOR2_X2 U1941 ( .A(n6529), .B(n255), .ZN(n1880) );
  OAI22_X2 U1942 ( .A1(n3954), .A2(n3368), .B1(n3953), .B2(n3952), .ZN(n3955)
         );
  NAND2_X2 U1943 ( .A1(n3538), .A2(a[15]), .ZN(n3954) );
  INV_X1 U1944 ( .A(n3482), .ZN(n3913) );
  NAND2_X2 U1945 ( .A1(n3202), .A2(n3082), .ZN(n780) );
  NOR2_X2 U1947 ( .A1(n4382), .A2(n2296), .ZN(n3015) );
  NAND3_X1 U1948 ( .A1(n314), .A2(n1190), .A3(n5427), .ZN(n5437) );
  NOR2_X1 U1949 ( .A1(n1599), .A2(n4582), .ZN(n1598) );
  NAND2_X2 U1950 ( .A1(n649), .A2(n650), .ZN(n652) );
  INV_X2 U1951 ( .A(n1571), .ZN(n649) );
  INV_X1 U1954 ( .A(n2824), .ZN(n654) );
  INV_X1 U1955 ( .A(n4671), .ZN(n2824) );
  NAND2_X1 U1956 ( .A1(n4216), .A2(b[6]), .ZN(n657) );
  NAND2_X1 U1957 ( .A1(n4217), .A2(n1324), .ZN(n658) );
  BUF_X4 U1960 ( .A(n2093), .Z(n1105) );
  NAND2_X1 U1963 ( .A1(n1698), .A2(n5330), .ZN(n661) );
  INV_X2 U1964 ( .A(n1698), .ZN(n659) );
  NAND2_X1 U1968 ( .A1(n1785), .A2(n4865), .ZN(n668) );
  NOR2_X2 U1974 ( .A1(n3431), .A2(b[7]), .ZN(n1554) );
  INV_X1 U1979 ( .A(n4633), .ZN(n675) );
  NAND2_X2 U1980 ( .A1(n1002), .A2(n6325), .ZN(n3625) );
  AOI22_X1 U1981 ( .A1(n4754), .A2(n4753), .B1(b[4]), .B2(n4752), .ZN(n3278)
         );
  NAND2_X1 U1982 ( .A1(n4308), .A2(n4244), .ZN(n678) );
  NAND2_X2 U1984 ( .A1(n3670), .A2(n2879), .ZN(n679) );
  NAND2_X1 U1986 ( .A1(n5077), .A2(b[0]), .ZN(n1741) );
  NAND2_X1 U1988 ( .A1(n1351), .A2(n5870), .ZN(n682) );
  NAND2_X2 U1989 ( .A1(n683), .A2(n682), .ZN(\d[39]_BAR ) );
  INV_X1 U1990 ( .A(n5870), .ZN(n681) );
  NAND2_X2 U1992 ( .A1(n5043), .A2(n5044), .ZN(n687) );
  NAND2_X2 U1993 ( .A1(n686), .A2(n687), .ZN(n3530) );
  NAND2_X1 U1996 ( .A1(n5610), .A2(n5869), .ZN(n5870) );
  NAND2_X1 U1997 ( .A1(n4871), .A2(n4968), .ZN(n691) );
  XNOR2_X2 U2002 ( .A(n4837), .B(n1215), .ZN(n1230) );
  NAND2_X4 U2009 ( .A1(a[5]), .A2(a[6]), .ZN(n702) );
  INV_X4 U2010 ( .A(a[5]), .ZN(n700) );
  INV_X8 U2011 ( .A(a[6]), .ZN(n701) );
  NAND2_X2 U2013 ( .A1(n3259), .A2(n3258), .ZN(n705) );
  NAND2_X4 U2015 ( .A1(n706), .A2(n705), .ZN(n5041) );
  INV_X2 U2016 ( .A(n3259), .ZN(n703) );
  NAND2_X2 U2018 ( .A1(n5041), .A2(b[21]), .ZN(n3587) );
  NAND2_X1 U2019 ( .A1(n1937), .A2(n4684), .ZN(n707) );
  NOR2_X1 U2021 ( .A1(n2578), .A2(n2588), .ZN(n5745) );
  INV_X1 U2022 ( .A(n2588), .ZN(n2516) );
  NOR2_X1 U2027 ( .A1(n1002), .A2(n5768), .ZN(n5769) );
  INV_X4 U2028 ( .A(n4909), .ZN(n1898) );
  NOR2_X2 U2029 ( .A1(n3680), .A2(n4909), .ZN(n1986) );
  NOR2_X4 U2030 ( .A1(n1134), .A2(n1133), .ZN(n3452) );
  OAI21_X2 U2032 ( .B1(n4038), .B2(n4037), .A(n3594), .ZN(n712) );
  NAND3_X1 U2033 ( .A1(n2368), .A2(n3060), .A3(n4470), .ZN(n2367) );
  NAND2_X1 U2034 ( .A1(n4961), .A2(n4962), .ZN(n714) );
  NAND2_X2 U2035 ( .A1(n4964), .A2(n713), .ZN(n715) );
  NAND2_X2 U2036 ( .A1(n714), .A2(n715), .ZN(n2576) );
  INV_X2 U2037 ( .A(n4962), .ZN(n713) );
  NAND2_X1 U2038 ( .A1(n2576), .A2(n6511), .ZN(n2883) );
  NAND2_X1 U2039 ( .A1(n4339), .A2(n6609), .ZN(n2180) );
  NAND2_X1 U2041 ( .A1(n5288), .A2(n5289), .ZN(n719) );
  NAND2_X2 U2042 ( .A1(n6152), .A2(n6150), .ZN(n720) );
  NAND2_X2 U2043 ( .A1(n719), .A2(n720), .ZN(n5238) );
  NAND2_X1 U2046 ( .A1(n1877), .A2(n41), .ZN(n723) );
  NAND2_X2 U2047 ( .A1(n721), .A2(n722), .ZN(n724) );
  NAND2_X2 U2048 ( .A1(n723), .A2(n724), .ZN(n5288) );
  INV_X2 U2049 ( .A(n1877), .ZN(n721) );
  OAI22_X2 U2051 ( .A1(n4999), .A2(b[12]), .B1(n3056), .B2(n3617), .ZN(n1564)
         );
  AOI22_X1 U2053 ( .A1(n5424), .A2(n6515), .B1(n1193), .B2(n3020), .ZN(n2408)
         );
  NAND2_X2 U2054 ( .A1(n2510), .A2(n2603), .ZN(n3907) );
  NAND2_X1 U2055 ( .A1(n3191), .A2(n3192), .ZN(n727) );
  NAND2_X2 U2056 ( .A1(n725), .A2(n5563), .ZN(n728) );
  INV_X2 U2058 ( .A(n3192), .ZN(n725) );
  INV_X1 U2061 ( .A(n5562), .ZN(n729) );
  INV_X4 U2062 ( .A(n4952), .ZN(n2303) );
  INV_X4 U2063 ( .A(n5014), .ZN(n1284) );
  NAND2_X4 U2064 ( .A1(n1066), .A2(n733), .ZN(n735) );
  NAND2_X4 U2065 ( .A1(n734), .A2(n735), .ZN(n3573) );
  INV_X8 U2066 ( .A(a[4]), .ZN(n733) );
  INV_X4 U2068 ( .A(n3573), .ZN(n1524) );
  NAND2_X1 U2069 ( .A1(n5315), .A2(n3371), .ZN(n736) );
  NAND2_X1 U2071 ( .A1(n2930), .A2(n4575), .ZN(n739) );
  NAND3_X2 U2074 ( .A1(n3838), .A2(n3764), .A3(n4271), .ZN(n3462) );
  NAND2_X2 U2075 ( .A1(n3834), .A2(n1287), .ZN(n3764) );
  NOR2_X4 U2076 ( .A1(n275), .A2(n3266), .ZN(n3264) );
  NAND2_X1 U2077 ( .A1(n2846), .A2(n5354), .ZN(n742) );
  NAND2_X2 U2078 ( .A1(n740), .A2(n741), .ZN(n743) );
  NAND2_X2 U2079 ( .A1(n742), .A2(n743), .ZN(n5330) );
  INV_X2 U2080 ( .A(n2846), .ZN(n740) );
  INV_X2 U2081 ( .A(n5354), .ZN(n741) );
  NAND2_X1 U2082 ( .A1(n2813), .A2(n2812), .ZN(n746) );
  INV_X1 U2084 ( .A(n2812), .ZN(n745) );
  INV_X1 U2085 ( .A(n2064), .ZN(n5354) );
  NAND2_X1 U2087 ( .A1(n473), .A2(n2899), .ZN(n1694) );
  OAI21_X1 U2088 ( .B1(n4058), .B2(n4057), .A(n4056), .ZN(n4067) );
  NAND2_X1 U2089 ( .A1(n5242), .A2(n748), .ZN(n749) );
  INV_X1 U2090 ( .A(n761), .ZN(n748) );
  NOR2_X1 U2091 ( .A1(n3509), .A2(n3346), .ZN(n751) );
  NOR2_X2 U2092 ( .A1(n3346), .A2(n3509), .ZN(n1281) );
  NOR2_X1 U2093 ( .A1(n1847), .A2(b[5]), .ZN(n3836) );
  NAND2_X1 U2094 ( .A1(n1847), .A2(n4614), .ZN(n4335) );
  NAND2_X1 U2096 ( .A1(n1847), .A2(n3020), .ZN(n2146) );
  INV_X8 U2097 ( .A(n2589), .ZN(n4483) );
  NOR2_X4 U2098 ( .A1(n2954), .A2(a[19]), .ZN(n2589) );
  NOR2_X1 U2100 ( .A1(n5670), .A2(n5671), .ZN(n5677) );
  NAND2_X1 U2101 ( .A1(n4650), .A2(n4651), .ZN(n1993) );
  NAND2_X2 U2102 ( .A1(n2163), .A2(n4488), .ZN(n4642) );
  NAND2_X1 U2103 ( .A1(n2324), .A2(n2719), .ZN(n756) );
  NAND2_X2 U2105 ( .A1(n1727), .A2(n4854), .ZN(n4862) );
  NAND2_X2 U2106 ( .A1(n4855), .A2(n4862), .ZN(n4856) );
  INV_X4 U2108 ( .A(n1378), .ZN(n759) );
  NOR2_X4 U2109 ( .A1(n937), .A2(a[17]), .ZN(n760) );
  INV_X4 U2113 ( .A(n3403), .ZN(n833) );
  AOI22_X1 U2114 ( .A1(n4705), .A2(b[8]), .B1(n3342), .B2(n998), .ZN(n1874) );
  INV_X1 U2115 ( .A(n2658), .ZN(n2882) );
  NAND2_X1 U2117 ( .A1(n3930), .A2(n3932), .ZN(n764) );
  INV_X1 U2121 ( .A(n3932), .ZN(n763) );
  NAND2_X1 U2122 ( .A1(n1593), .A2(n3936), .ZN(n769) );
  INV_X2 U2125 ( .A(n1593), .ZN(n767) );
  AOI22_X1 U2126 ( .A1(n3896), .A2(n3895), .B1(n967), .B2(n1010), .ZN(n3932)
         );
  NAND2_X2 U2128 ( .A1(n772), .A2(n773), .ZN(n775) );
  INV_X1 U2131 ( .A(n2087), .ZN(n4649) );
  INV_X1 U2132 ( .A(n4737), .ZN(n2311) );
  INV_X2 U2134 ( .A(n2773), .ZN(n777) );
  INV_X1 U2136 ( .A(n4538), .ZN(n3713) );
  NAND2_X2 U2137 ( .A1(n324), .A2(n1581), .ZN(n807) );
  BUF_X4 U2138 ( .A(n3082), .Z(n781) );
  NAND3_X2 U2141 ( .A1(n4159), .A2(n4559), .A3(a[0]), .ZN(n2097) );
  AOI22_X1 U2142 ( .A1(n4159), .A2(a[0]), .B1(n4219), .B2(n3465), .ZN(n4161)
         );
  NAND2_X2 U2143 ( .A1(n2246), .A2(n2245), .ZN(n782) );
  NAND3_X1 U2145 ( .A1(n1039), .A2(n2322), .A3(n3928), .ZN(n2444) );
  NAND2_X1 U2146 ( .A1(n2074), .A2(n2073), .ZN(n785) );
  INV_X2 U2150 ( .A(n2073), .ZN(n784) );
  NAND2_X2 U2151 ( .A1(n3580), .A2(n2083), .ZN(n787) );
  NAND2_X2 U2153 ( .A1(n2932), .A2(n3342), .ZN(n1983) );
  NAND2_X2 U2155 ( .A1(n3528), .A2(n3529), .ZN(n790) );
  AOI21_X1 U2156 ( .B1(n3522), .B2(n3521), .A(n3523), .ZN(n1637) );
  INV_X4 U2161 ( .A(n1836), .ZN(n1201) );
  OAI21_X1 U2165 ( .B1(n3607), .B2(n3598), .A(n3284), .ZN(n2839) );
  NAND2_X2 U2172 ( .A1(n3013), .A2(n800), .ZN(n802) );
  INV_X4 U2175 ( .A(n4652), .ZN(n800) );
  NAND2_X1 U2177 ( .A1(n1943), .A2(n6200), .ZN(n803) );
  NAND2_X2 U2178 ( .A1(n804), .A2(n803), .ZN(n1942) );
  INV_X1 U2179 ( .A(n3480), .ZN(n1943) );
  INV_X1 U2181 ( .A(n4435), .ZN(n2159) );
  NAND2_X1 U2182 ( .A1(n1299), .A2(n4900), .ZN(n1300) );
  NAND2_X2 U2186 ( .A1(n5090), .A2(n5089), .ZN(n2799) );
  AOI22_X1 U2187 ( .A1(n2510), .A2(n6569), .B1(n2382), .B2(b[1]), .ZN(n3957)
         );
  AOI22_X1 U2188 ( .A1(n4145), .A2(n4144), .B1(n4143), .B2(n4142), .ZN(n5658)
         );
  NAND2_X2 U2192 ( .A1(n2743), .A2(n1059), .ZN(n3224) );
  NAND2_X2 U2196 ( .A1(n815), .A2(n816), .ZN(n964) );
  NAND2_X1 U2198 ( .A1(n328), .A2(n4942), .ZN(n1113) );
  OAI21_X1 U2199 ( .B1(n5276), .B2(n5275), .A(n2562), .ZN(n2559) );
  NOR3_X1 U2200 ( .A1(n5276), .A2(n5275), .A3(n2562), .ZN(n2561) );
  NOR2_X2 U2207 ( .A1(n5665), .A2(n4152), .ZN(n4151) );
  NOR2_X1 U2208 ( .A1(n3573), .A2(n3905), .ZN(n2307) );
  NAND2_X1 U2210 ( .A1(n6456), .A2(n3131), .ZN(n1322) );
  INV_X4 U2211 ( .A(n5212), .ZN(n821) );
  NAND2_X2 U2213 ( .A1(n825), .A2(n826), .ZN(n828) );
  NAND2_X2 U2214 ( .A1(n827), .A2(n6514), .ZN(n5090) );
  NAND2_X2 U2217 ( .A1(n980), .A2(n979), .ZN(n978) );
  NAND2_X2 U2220 ( .A1(n831), .A2(n832), .ZN(n5060) );
  INV_X1 U2221 ( .A(n5117), .ZN(n830) );
  NAND2_X1 U2223 ( .A1(n2544), .A2(n4000), .ZN(n838) );
  NAND2_X2 U2224 ( .A1(n836), .A2(n837), .ZN(n839) );
  INV_X1 U2227 ( .A(n4000), .ZN(n837) );
  NAND2_X4 U2229 ( .A1(a[8]), .A2(a[7]), .ZN(n845) );
  NAND2_X4 U2230 ( .A1(n843), .A2(n844), .ZN(n846) );
  NAND2_X4 U2231 ( .A1(n846), .A2(n845), .ZN(n3395) );
  INV_X4 U2232 ( .A(a[8]), .ZN(n843) );
  INV_X8 U2233 ( .A(a[7]), .ZN(n844) );
  NAND2_X1 U2236 ( .A1(n4387), .A2(n4388), .ZN(n1141) );
  NAND2_X1 U2241 ( .A1(n4175), .A2(n1626), .ZN(n4197) );
  NAND3_X1 U2242 ( .A1(n1783), .A2(n2076), .A3(n2360), .ZN(n1782) );
  NAND2_X1 U2243 ( .A1(n5113), .A2(n2360), .ZN(n1781) );
  NAND2_X1 U2244 ( .A1(n2360), .A2(n2354), .ZN(n1780) );
  INV_X1 U2251 ( .A(n5777), .ZN(n5765) );
  NOR2_X2 U2252 ( .A1(n5764), .A2(n5772), .ZN(n5777) );
  NAND2_X1 U2253 ( .A1(n2113), .A2(n4279), .ZN(n855) );
  NAND2_X2 U2254 ( .A1(n853), .A2(n854), .ZN(n856) );
  INV_X2 U2256 ( .A(n2113), .ZN(n853) );
  INV_X1 U2257 ( .A(n4279), .ZN(n854) );
  NAND3_X1 U2260 ( .A1(n3325), .A2(n5176), .A3(n2401), .ZN(n1630) );
  NAND2_X4 U2261 ( .A1(a[23]), .A2(b[2]), .ZN(n4724) );
  NAND2_X2 U2262 ( .A1(n857), .A2(n6504), .ZN(n860) );
  NAND2_X1 U2264 ( .A1(n2239), .A2(n4275), .ZN(n863) );
  INV_X2 U2267 ( .A(n2239), .ZN(n861) );
  INV_X1 U2268 ( .A(n4275), .ZN(n862) );
  NAND2_X4 U2269 ( .A1(n6608), .A2(n4924), .ZN(n4796) );
  INV_X4 U2272 ( .A(n3463), .ZN(n2140) );
  NAND2_X1 U2273 ( .A1(n3838), .A2(n3764), .ZN(n4272) );
  NOR2_X1 U2274 ( .A1(n3806), .A2(n6215), .ZN(n3807) );
  NAND2_X2 U2276 ( .A1(n866), .A2(n867), .ZN(n869) );
  INV_X4 U2279 ( .A(n2291), .ZN(n870) );
  INV_X4 U2283 ( .A(n1540), .ZN(n873) );
  NAND2_X2 U2286 ( .A1(n877), .A2(n4906), .ZN(n880) );
  INV_X2 U2288 ( .A(n3219), .ZN(n877) );
  NAND3_X1 U2290 ( .A1(n3291), .A2(n3290), .A3(n3268), .ZN(n1858) );
  NAND2_X2 U2292 ( .A1(n1903), .A2(n1905), .ZN(n881) );
  NOR2_X1 U2293 ( .A1(n3854), .A2(n1000), .ZN(n2748) );
  NAND2_X1 U2296 ( .A1(n2167), .A2(n2168), .ZN(n1247) );
  NAND2_X4 U2297 ( .A1(n2683), .A2(n2682), .ZN(n4765) );
  NAND2_X2 U2299 ( .A1(n388), .A2(n6519), .ZN(n882) );
  NAND2_X1 U2300 ( .A1(n2966), .A2(n971), .ZN(n885) );
  NAND2_X1 U2304 ( .A1(n2205), .A2(n5246), .ZN(n889) );
  INV_X2 U2307 ( .A(n2205), .ZN(n887) );
  NOR2_X1 U2309 ( .A1(n3867), .A2(n3868), .ZN(n2308) );
  AOI22_X2 U2310 ( .A1(n1942), .A2(n1112), .B1(n1941), .B2(n5039), .ZN(n891)
         );
  NAND2_X4 U2320 ( .A1(n1224), .A2(n1223), .ZN(n4908) );
  INV_X1 U2321 ( .A(n283), .ZN(n2578) );
  AOI22_X2 U2322 ( .A1(n2084), .A2(n3561), .B1(n2085), .B2(n6655), .ZN(n2083)
         );
  INV_X4 U2323 ( .A(n4382), .ZN(n2543) );
  NAND2_X2 U2324 ( .A1(n5699), .A2(n3365), .ZN(n903) );
  INV_X1 U2330 ( .A(n2508), .ZN(n1124) );
  NAND2_X1 U2331 ( .A1(n758), .A2(b[14]), .ZN(n2077) );
  NAND2_X1 U2335 ( .A1(n2369), .A2(n4872), .ZN(n914) );
  NAND2_X2 U2336 ( .A1(n912), .A2(n913), .ZN(n915) );
  NAND2_X2 U2337 ( .A1(n915), .A2(n914), .ZN(n2410) );
  INV_X2 U2338 ( .A(n2369), .ZN(n912) );
  INV_X4 U2340 ( .A(n1025), .ZN(n916) );
  NAND2_X4 U2343 ( .A1(a[13]), .A2(a[14]), .ZN(n919) );
  NAND2_X4 U2344 ( .A1(n917), .A2(n918), .ZN(n920) );
  NAND2_X4 U2345 ( .A1(n920), .A2(n919), .ZN(n5197) );
  INV_X4 U2346 ( .A(a[13]), .ZN(n917) );
  INV_X8 U2347 ( .A(a[14]), .ZN(n918) );
  NOR2_X1 U2348 ( .A1(n4504), .A2(n3465), .ZN(n923) );
  OAI21_X1 U2350 ( .B1(n6525), .B2(n5884), .A(n5883), .ZN(n5886) );
  NAND2_X2 U2351 ( .A1(n925), .A2(n926), .ZN(n928) );
  NAND2_X2 U2352 ( .A1(n927), .A2(n928), .ZN(\d[38]_BAR ) );
  NAND2_X2 U2354 ( .A1(n930), .A2(n931), .ZN(n2004) );
  NAND2_X2 U2357 ( .A1(n932), .A2(n531), .ZN(n934) );
  NAND2_X4 U2359 ( .A1(a[16]), .A2(a[15]), .ZN(n937) );
  NOR2_X1 U2361 ( .A1(n5875), .A2(n5571), .ZN(n5373) );
  NAND2_X2 U2362 ( .A1(n2323), .A2(n2720), .ZN(n941) );
  NAND2_X1 U2364 ( .A1(n4509), .A2(n1935), .ZN(n944) );
  XNOR2_X1 U2369 ( .A(a[11]), .B(b[15]), .ZN(n4593) );
  XNOR2_X1 U2371 ( .A(a[9]), .B(b[21]), .ZN(n4770) );
  INV_X1 U2372 ( .A(n4726), .ZN(n4681) );
  NAND2_X1 U2373 ( .A1(b[5]), .A2(a[23]), .ZN(n4749) );
  INV_X1 U2378 ( .A(n4611), .ZN(n3292) );
  INV_X1 U2379 ( .A(n4880), .ZN(n1864) );
  NAND2_X2 U2381 ( .A1(n1524), .A2(n2709), .ZN(n3095) );
  NAND2_X1 U2382 ( .A1(n568), .A2(n5293), .ZN(n2017) );
  XNOR2_X1 U2385 ( .A(a[23]), .B(b[13]), .ZN(n5189) );
  NOR2_X1 U2388 ( .A1(n5190), .A2(n5189), .ZN(n5191) );
  NAND2_X1 U2391 ( .A1(n47), .A2(b[4]), .ZN(n1887) );
  NAND2_X1 U2392 ( .A1(a[8]), .A2(b[3]), .ZN(n3539) );
  NAND2_X1 U2393 ( .A1(n2753), .A2(n2752), .ZN(n2750) );
  NAND2_X1 U2394 ( .A1(n6035), .A2(n5293), .ZN(n3515) );
  NAND2_X1 U2397 ( .A1(n4365), .A2(b[0]), .ZN(n3794) );
  NOR2_X1 U2398 ( .A1(n3728), .A2(b[1]), .ZN(n1823) );
  NAND2_X1 U2400 ( .A1(n4746), .A2(n4598), .ZN(n1210) );
  NOR2_X1 U2401 ( .A1(b[0]), .A2(n4600), .ZN(n1919) );
  NAND2_X1 U2404 ( .A1(n5563), .A2(n5562), .ZN(n5559) );
  INV_X1 U2405 ( .A(n5958), .ZN(n5959) );
  NAND2_X1 U2407 ( .A1(n6198), .A2(n2573), .ZN(n1663) );
  NOR2_X1 U2410 ( .A1(n5774), .A2(n5771), .ZN(n5766) );
  NAND2_X1 U2411 ( .A1(n6097), .A2(n4133), .ZN(n5652) );
  XNOR2_X2 U2418 ( .A(a[5]), .B(b[1]), .ZN(n950) );
  AND3_X1 U2420 ( .A1(n4009), .A2(n3202), .A3(n3082), .ZN(n952) );
  NAND2_X2 U2422 ( .A1(n1132), .A2(n4729), .ZN(n1146) );
  OR2_X4 U2423 ( .A1(n5149), .A2(n5150), .ZN(n954) );
  INV_X1 U2429 ( .A(n5011), .ZN(n4958) );
  INV_X1 U2430 ( .A(n5717), .ZN(n1021) );
  INV_X1 U2431 ( .A(n5177), .ZN(n3325) );
  XOR2_X2 U2434 ( .A(b[7]), .B(a[1]), .Z(n961) );
  INV_X1 U2437 ( .A(n3922), .ZN(n2845) );
  OR2_X4 U2439 ( .A1(n2345), .A2(n5501), .ZN(n966) );
  AND2_X4 U2440 ( .A1(n1514), .A2(n3890), .ZN(n967) );
  OR2_X4 U2442 ( .A1(n5472), .A2(n5951), .ZN(n970) );
  AND2_X2 U2445 ( .A1(n4842), .A2(n4841), .ZN(n973) );
  OAI21_X1 U2446 ( .B1(n975), .B2(b[5]), .A(n974), .ZN(n4186) );
  NAND2_X1 U2447 ( .A1(n4504), .A2(b[5]), .ZN(n974) );
  NAND3_X1 U2449 ( .A1(n3117), .A2(n6062), .A3(n1902), .ZN(n3611) );
  NOR2_X1 U2450 ( .A1(n472), .A2(b[12]), .ZN(n3555) );
  INV_X2 U2451 ( .A(a[8]), .ZN(n980) );
  OAI21_X1 U2452 ( .B1(n975), .B2(b[11]), .A(n983), .ZN(n3853) );
  NAND2_X1 U2453 ( .A1(b[11]), .A2(n4504), .ZN(n983) );
  OR2_X2 U2454 ( .A1(n5899), .A2(n984), .ZN(n2055) );
  INV_X1 U2459 ( .A(n4938), .ZN(n2659) );
  NAND2_X1 U2460 ( .A1(n4671), .A2(n1119), .ZN(n2230) );
  AND2_X4 U2464 ( .A1(n47), .A2(b[10]), .ZN(n992) );
  INV_X1 U2465 ( .A(n4315), .ZN(n4006) );
  AND2_X4 U2466 ( .A1(n6622), .A2(n4738), .ZN(n994) );
  NAND2_X1 U2469 ( .A1(n1545), .A2(n3640), .ZN(n1471) );
  XNOR2_X2 U2470 ( .A(a[10]), .B(a[9]), .ZN(n999) );
  XNOR2_X2 U2471 ( .A(a[10]), .B(a[9]), .ZN(n1000) );
  INV_X2 U2472 ( .A(n6021), .ZN(n6022) );
  NAND2_X2 U2473 ( .A1(n3476), .A2(n6016), .ZN(n6017) );
  INV_X2 U2474 ( .A(n5778), .ZN(n5773) );
  INV_X2 U2475 ( .A(n5827), .ZN(n5816) );
  INV_X4 U2478 ( .A(n1068), .ZN(n1651) );
  INV_X2 U2479 ( .A(n3525), .ZN(n1641) );
  AOI22_X2 U2480 ( .A1(n5489), .A2(n5486), .B1(n5485), .B2(n5487), .ZN(n5574)
         );
  XNOR2_X2 U2483 ( .A(n1315), .B(n3705), .ZN(n5680) );
  INV_X4 U2484 ( .A(n5307), .ZN(n1001) );
  NAND2_X1 U2485 ( .A1(n5937), .A2(n5936), .ZN(n6075) );
  NAND2_X1 U2486 ( .A1(n5690), .A2(n1008), .ZN(n5692) );
  XNOR2_X1 U2488 ( .A(n5912), .B(n5911), .ZN(n5935) );
  INV_X2 U2489 ( .A(n5502), .ZN(n5463) );
  NOR2_X1 U2490 ( .A1(n4201), .A2(n5670), .ZN(n4200) );
  INV_X4 U2491 ( .A(n4072), .ZN(n2636) );
  INV_X2 U2492 ( .A(n4954), .ZN(n4955) );
  INV_X2 U2493 ( .A(n4953), .ZN(n4957) );
  NAND2_X1 U2494 ( .A1(n5510), .A2(n5480), .ZN(n5482) );
  NOR2_X1 U2495 ( .A1(n5510), .A2(n5480), .ZN(n5481) );
  NAND2_X1 U2496 ( .A1(n4378), .A2(n4379), .ZN(n4381) );
  INV_X2 U2497 ( .A(n5908), .ZN(n5909) );
  INV_X2 U2498 ( .A(n5349), .ZN(n5350) );
  OR2_X2 U2499 ( .A1(n967), .A2(n1010), .ZN(n3896) );
  NAND2_X2 U2502 ( .A1(n5224), .A2(n3011), .ZN(n5296) );
  NAND2_X1 U2503 ( .A1(n3272), .A2(n3271), .ZN(n3270) );
  NOR2_X1 U2509 ( .A1(n2213), .A2(n2212), .ZN(n2211) );
  NAND2_X2 U2510 ( .A1(n3330), .A2(n3329), .ZN(n4507) );
  INV_X1 U2511 ( .A(n4617), .ZN(n4618) );
  OR2_X2 U2512 ( .A1(n4835), .A2(n4834), .ZN(n1251) );
  INV_X2 U2513 ( .A(n3610), .ZN(n3156) );
  XOR2_X2 U2518 ( .A(b[8]), .B(a[19]), .Z(n4688) );
  XOR2_X2 U2519 ( .A(b[17]), .B(a[13]), .Z(n4775) );
  INV_X2 U2521 ( .A(b[6]), .ZN(n4011) );
  XNOR2_X1 U2522 ( .A(b[10]), .B(a[1]), .ZN(n4221) );
  XOR2_X2 U2525 ( .A(a[15]), .B(b[2]), .Z(n3865) );
  XNOR2_X1 U2530 ( .A(a[1]), .B(b[3]), .ZN(n4132) );
  XOR2_X2 U2531 ( .A(a[11]), .B(b[11]), .Z(n4326) );
  INV_X4 U2532 ( .A(b[7]), .ZN(n3465) );
  XOR2_X2 U2534 ( .A(b[18]), .B(a[11]), .Z(n3261) );
  XOR2_X2 U2535 ( .A(a[11]), .B(b[2]), .Z(n3830) );
  INV_X1 U2537 ( .A(n6070), .ZN(n5872) );
  AND2_X2 U2539 ( .A1(n5861), .A2(n3719), .ZN(n3718) );
  NOR2_X1 U2542 ( .A1(n5750), .A2(n5758), .ZN(n5752) );
  INV_X2 U2543 ( .A(n5389), .ZN(n3392) );
  INV_X2 U2546 ( .A(n5713), .ZN(n5703) );
  AOI21_X1 U2547 ( .B1(n5706), .B2(n5711), .A(n5713), .ZN(n5709) );
  NOR2_X2 U2549 ( .A1(n5698), .A2(n5697), .ZN(n5702) );
  INV_X2 U2550 ( .A(n5091), .ZN(n2420) );
  INV_X4 U2551 ( .A(n3474), .ZN(n1400) );
  INV_X2 U2553 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U2554 ( .A1(n1020), .A2(n6075), .ZN(n6076) );
  INV_X2 U2555 ( .A(n6074), .ZN(n1020) );
  NAND2_X2 U2557 ( .A1(n6064), .A2(n6065), .ZN(n6074) );
  NAND2_X2 U2560 ( .A1(n5934), .A2(n5935), .ZN(n6065) );
  INV_X1 U2561 ( .A(n5935), .ZN(n5936) );
  INV_X1 U2562 ( .A(n5934), .ZN(n5937) );
  NOR2_X1 U2563 ( .A1(n6112), .A2(n6117), .ZN(n6110) );
  INV_X4 U2564 ( .A(n3615), .ZN(n1003) );
  NAND2_X2 U2566 ( .A1(n2231), .A2(n2230), .ZN(n4733) );
  OAI21_X1 U2567 ( .B1(n5891), .B2(n5890), .A(n5889), .ZN(n5934) );
  INV_X2 U2568 ( .A(n2880), .ZN(n4963) );
  INV_X2 U2569 ( .A(n5133), .ZN(n1031) );
  NAND2_X4 U2570 ( .A1(n1161), .A2(n1160), .ZN(n2937) );
  OAI21_X1 U2571 ( .B1(n5537), .B2(n5536), .A(n5535), .ZN(n5538) );
  NAND2_X1 U2572 ( .A1(n5893), .A2(n5892), .ZN(n5940) );
  INV_X2 U2573 ( .A(n4738), .ZN(n2833) );
  INV_X2 U2575 ( .A(n4459), .ZN(n4460) );
  INV_X4 U2576 ( .A(n4669), .ZN(n1005) );
  INV_X1 U2577 ( .A(n6027), .ZN(n6028) );
  INV_X4 U2578 ( .A(n1036), .ZN(n1007) );
  INV_X2 U2579 ( .A(n4571), .ZN(n1977) );
  INV_X2 U2580 ( .A(n5509), .ZN(n5480) );
  XNOR2_X1 U2581 ( .A(n1681), .B(n1680), .ZN(n5412) );
  INV_X2 U2582 ( .A(n4859), .ZN(n1250) );
  INV_X1 U2583 ( .A(n5438), .ZN(n5428) );
  INV_X2 U2585 ( .A(n5175), .ZN(n1042) );
  NOR2_X2 U2586 ( .A1(n6032), .A2(n5950), .ZN(n5955) );
  XNOR2_X1 U2587 ( .A(n5517), .B(n5516), .ZN(n1681) );
  OAI21_X1 U2588 ( .B1(n2399), .B2(n1255), .A(n1062), .ZN(n1253) );
  INV_X2 U2589 ( .A(n4720), .ZN(n4663) );
  NAND2_X1 U2590 ( .A1(n2820), .A2(n2819), .ZN(n5441) );
  INV_X1 U2594 ( .A(n6032), .ZN(n6037) );
  INV_X2 U2595 ( .A(n4622), .ZN(n4623) );
  NAND2_X1 U2596 ( .A1(n5340), .A2(n2932), .ZN(n5449) );
  INV_X2 U2598 ( .A(n2549), .ZN(n4807) );
  INV_X4 U2599 ( .A(n3894), .ZN(n1010) );
  INV_X1 U2600 ( .A(n4141), .ZN(n4143) );
  NOR2_X2 U2602 ( .A1(n2594), .A2(n2593), .ZN(n1801) );
  MUX2_X2 U2603 ( .A(n2514), .B(n5526), .S(n5105), .Z(n5527) );
  NAND2_X1 U2609 ( .A1(n2097), .A2(n2096), .ZN(n2095) );
  INV_X2 U2610 ( .A(n4031), .ZN(n1057) );
  NAND2_X1 U2613 ( .A1(n4618), .A2(n4619), .ZN(n2466) );
  NAND2_X1 U2614 ( .A1(n2932), .A2(n2569), .ZN(n2568) );
  NAND2_X2 U2615 ( .A1(n1542), .A2(a[0]), .ZN(n1539) );
  INV_X1 U2616 ( .A(n5422), .ZN(n3547) );
  MUX2_X2 U2617 ( .A(n5531), .B(n5530), .S(b[19]), .Z(n5532) );
  NAND2_X2 U2619 ( .A1(n6038), .A2(n5953), .ZN(n5954) );
  INV_X1 U2620 ( .A(n5020), .ZN(n5022) );
  INV_X4 U2621 ( .A(n4767), .ZN(n5424) );
  AOI21_X1 U2623 ( .B1(b[9]), .B2(b[8]), .A(n5151), .ZN(n5080) );
  AND2_X1 U2624 ( .A1(a[19]), .A2(n984), .ZN(n2749) );
  INV_X8 U2625 ( .A(n4543), .ZN(n1012) );
  INV_X2 U2626 ( .A(n4873), .ZN(n1063) );
  INV_X2 U2629 ( .A(b[5]), .ZN(n1884) );
  INV_X2 U2630 ( .A(b[7]), .ZN(n4687) );
  INV_X4 U2632 ( .A(a[9]), .ZN(n3058) );
  XOR2_X2 U2634 ( .A(b[12]), .B(a[13]), .Z(n4529) );
  XOR2_X2 U2635 ( .A(a[15]), .B(b[10]), .Z(n4530) );
  XOR2_X2 U2636 ( .A(a[11]), .B(b[14]), .Z(n4558) );
  XOR2_X2 U2637 ( .A(a[5]), .B(b[17]), .Z(n4317) );
  XOR2_X2 U2639 ( .A(a[5]), .B(b[10]), .Z(n3785) );
  NAND2_X2 U2641 ( .A1(a[23]), .A2(b[10]), .ZN(n5166) );
  XOR2_X2 U2642 ( .A(b[7]), .B(a[7]), .Z(n3803) );
  XOR2_X1 U2643 ( .A(b[8]), .B(a[5]), .Z(n3840) );
  XOR2_X2 U2644 ( .A(a[11]), .B(b[9]), .Z(n4025) );
  XNOR2_X1 U2645 ( .A(b[5]), .B(a[1]), .ZN(n4111) );
  INV_X2 U2647 ( .A(n1327), .ZN(n5387) );
  INV_X2 U2649 ( .A(n6080), .ZN(n6083) );
  INV_X2 U2650 ( .A(n6009), .ZN(n6011) );
  INV_X2 U2652 ( .A(n5590), .ZN(n5588) );
  OR2_X2 U2653 ( .A1(n6016), .A2(n3724), .ZN(n3725) );
  INV_X2 U2654 ( .A(n6016), .ZN(n6014) );
  INV_X4 U2655 ( .A(n5928), .ZN(n1013) );
  INV_X2 U2656 ( .A(n5980), .ZN(n5991) );
  AND2_X2 U2657 ( .A1(n2864), .A2(n5855), .ZN(n3099) );
  NAND2_X1 U2658 ( .A1(n5732), .A2(n5731), .ZN(n5739) );
  NOR2_X1 U2661 ( .A1(n5931), .A2(n5932), .ZN(n2863) );
  AOI22_X1 U2662 ( .A1(n5752), .A2(n5751), .B1(n5753), .B2(n5750), .ZN(n5755)
         );
  INV_X2 U2665 ( .A(n1314), .ZN(n5877) );
  NAND2_X2 U2666 ( .A1(n2976), .A2(n5852), .ZN(n5855) );
  INV_X2 U2667 ( .A(n5829), .ZN(n5815) );
  INV_X2 U2670 ( .A(n5806), .ZN(n5807) );
  INV_X2 U2673 ( .A(n5760), .ZN(n5750) );
  XNOR2_X1 U2674 ( .A(n5709), .B(n5708), .ZN(\d[13]_BAR ) );
  NAND2_X2 U2675 ( .A1(n5703), .A2(n5711), .ZN(n5705) );
  INV_X2 U2676 ( .A(n5813), .ZN(n5821) );
  INV_X2 U2677 ( .A(n6084), .ZN(n6085) );
  INV_X2 U2680 ( .A(n5634), .ZN(n5635) );
  AOI22_X1 U2682 ( .A1(n5576), .A2(n5582), .B1(n5933), .B2(n5575), .ZN(n5577)
         );
  NOR2_X2 U2684 ( .A1(n3133), .A2(n1307), .ZN(n5713) );
  NAND2_X2 U2685 ( .A1(n3133), .A2(n1307), .ZN(n5711) );
  NOR2_X2 U2687 ( .A1(n6063), .A2(n5933), .ZN(n6078) );
  AND2_X2 U2688 ( .A1(n6063), .A2(n6064), .ZN(n6073) );
  INV_X2 U2689 ( .A(n5971), .ZN(n5972) );
  INV_X4 U2691 ( .A(n5324), .ZN(n1016) );
  INV_X1 U2692 ( .A(n5745), .ZN(n5726) );
  OAI21_X1 U2693 ( .B1(n5696), .B2(n5692), .A(n5691), .ZN(n5698) );
  INV_X2 U2694 ( .A(n5578), .ZN(n5581) );
  INV_X2 U2695 ( .A(n2243), .ZN(n3602) );
  INV_X2 U2696 ( .A(n5913), .ZN(n5994) );
  INV_X2 U2697 ( .A(n5772), .ZN(n5771) );
  NAND2_X2 U2698 ( .A1(n2299), .A2(n3619), .ZN(n1289) );
  INV_X4 U2699 ( .A(n3125), .ZN(n1017) );
  INV_X1 U2700 ( .A(n368), .ZN(n3383) );
  INV_X2 U2701 ( .A(n5215), .ZN(n5217) );
  INV_X2 U2702 ( .A(n4631), .ZN(n2666) );
  INV_X2 U2704 ( .A(n4642), .ZN(n1018) );
  INV_X2 U2705 ( .A(n5704), .ZN(n5706) );
  INV_X2 U2706 ( .A(n4079), .ZN(n2389) );
  OAI21_X1 U2708 ( .B1(n5563), .B2(n5562), .A(n5558), .ZN(n5560) );
  INV_X2 U2709 ( .A(n6129), .ZN(n6130) );
  OAI22_X1 U2710 ( .A1(n6128), .A2(n6127), .B1(n6126), .B2(n6125), .ZN(n6129)
         );
  INV_X2 U2712 ( .A(n5545), .ZN(n5543) );
  NAND2_X2 U2714 ( .A1(n5545), .A2(n5544), .ZN(n6064) );
  INV_X2 U2715 ( .A(n5544), .ZN(n5542) );
  AOI21_X1 U2716 ( .B1(n6118), .B2(n6117), .A(n6116), .ZN(n6127) );
  INV_X2 U2717 ( .A(n5032), .ZN(n1636) );
  NOR2_X1 U2718 ( .A1(n6110), .A2(n6051), .ZN(n6059) );
  NAND2_X2 U2719 ( .A1(n2881), .A2(n2882), .ZN(n2884) );
  INV_X4 U2720 ( .A(n5331), .ZN(n1023) );
  AND2_X2 U2722 ( .A1(n4006), .A2(n4007), .ZN(n2742) );
  INV_X4 U2726 ( .A(n3410), .ZN(n1024) );
  INV_X4 U2727 ( .A(n4900), .ZN(n1025) );
  INV_X1 U2728 ( .A(n6112), .ZN(n6116) );
  NAND2_X1 U2729 ( .A1(n6337), .A2(n69), .ZN(n5695) );
  XNOR2_X1 U2730 ( .A(n2984), .B(n5664), .ZN(n5669) );
  NOR2_X2 U2731 ( .A1(n4280), .A2(n4281), .ZN(n2286) );
  INV_X1 U2732 ( .A(n6115), .ZN(n6118) );
  INV_X2 U2733 ( .A(n5264), .ZN(n2497) );
  AOI21_X1 U2735 ( .B1(n6120), .B2(n6121), .A(n6119), .ZN(n6126) );
  INV_X2 U2737 ( .A(n4201), .ZN(n4202) );
  NOR2_X1 U2738 ( .A1(n6107), .A2(n6124), .ZN(n6113) );
  INV_X1 U2740 ( .A(n6051), .ZN(n6052) );
  INV_X4 U2741 ( .A(n4487), .ZN(n1027) );
  INV_X4 U2744 ( .A(n2805), .ZN(n1028) );
  INV_X2 U2745 ( .A(n5538), .ZN(n5890) );
  NAND2_X1 U2746 ( .A1(n6124), .A2(n6109), .ZN(n6115) );
  INV_X2 U2747 ( .A(n5433), .ZN(n5431) );
  INV_X2 U2749 ( .A(n5484), .ZN(n5487) );
  NAND2_X1 U2751 ( .A1(n6122), .A2(n6121), .ZN(n6109) );
  INV_X2 U2754 ( .A(n5551), .ZN(n5508) );
  NOR2_X1 U2755 ( .A1(n6122), .A2(n6121), .ZN(n6107) );
  INV_X4 U2756 ( .A(n1805), .ZN(n1032) );
  OAI21_X1 U2757 ( .B1(n6332), .B2(n5670), .A(n4197), .ZN(n4177) );
  NAND2_X2 U2758 ( .A1(n5352), .A2(n3660), .ZN(n2557) );
  MUX2_X2 U2760 ( .A(n6100), .B(n6099), .S(n6098), .Z(\d[3] ) );
  INV_X2 U2761 ( .A(n4468), .ZN(n4462) );
  NAND2_X2 U2762 ( .A1(n4461), .A2(n4460), .ZN(n4467) );
  NOR2_X1 U2763 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  INV_X2 U2764 ( .A(n5537), .ZN(n5404) );
  INV_X2 U2767 ( .A(n5941), .ZN(n5945) );
  INV_X2 U2768 ( .A(n5939), .ZN(n5943) );
  INV_X2 U2769 ( .A(n5511), .ZN(n5483) );
  INV_X2 U2770 ( .A(n5282), .ZN(n2663) );
  INV_X4 U2771 ( .A(n3987), .ZN(n1033) );
  INV_X2 U2773 ( .A(n3634), .ZN(n1034) );
  INV_X2 U2775 ( .A(n5460), .ZN(n5461) );
  NOR2_X1 U2777 ( .A1(n6103), .A2(n6102), .ZN(n6048) );
  INV_X2 U2778 ( .A(n5029), .ZN(n1035) );
  INV_X2 U2780 ( .A(n6097), .ZN(n4134) );
  INV_X2 U2781 ( .A(n5907), .ZN(n5910) );
  NAND2_X2 U2782 ( .A1(n1335), .A2(n1523), .ZN(n2888) );
  INV_X4 U2783 ( .A(n5285), .ZN(n5282) );
  INV_X4 U2784 ( .A(n5251), .ZN(n1036) );
  OAI21_X1 U2785 ( .B1(n5436), .B2(n5428), .A(n5437), .ZN(n5435) );
  NAND2_X2 U2786 ( .A1(n3112), .A2(n2703), .ZN(n3529) );
  NAND2_X1 U2787 ( .A1(n5517), .A2(n5516), .ZN(n1676) );
  AOI21_X1 U2789 ( .B1(n6037), .B2(n6041), .A(n6036), .ZN(n6103) );
  NAND2_X2 U2790 ( .A1(n3548), .A2(n3547), .ZN(n3766) );
  NAND2_X1 U2792 ( .A1(n4169), .A2(n4168), .ZN(n4170) );
  INV_X2 U2793 ( .A(n5494), .ZN(n5447) );
  INV_X2 U2794 ( .A(n5273), .ZN(n5271) );
  INV_X2 U2795 ( .A(n5523), .ZN(n5521) );
  INV_X2 U2796 ( .A(n5956), .ZN(n5961) );
  INV_X2 U2797 ( .A(n4785), .ZN(n4786) );
  INV_X2 U2798 ( .A(n4040), .ZN(n4041) );
  NAND2_X2 U2799 ( .A1(n1490), .A2(n1011), .ZN(n3751) );
  INV_X2 U2801 ( .A(n3017), .ZN(n3016) );
  INV_X4 U2803 ( .A(n4621), .ZN(n1040) );
  NOR2_X2 U2804 ( .A1(n4020), .A2(n4019), .ZN(n2992) );
  NAND2_X2 U2805 ( .A1(n1252), .A2(n1251), .ZN(n4859) );
  INV_X2 U2808 ( .A(n4055), .ZN(n4064) );
  NOR2_X1 U2811 ( .A1(n3797), .A2(n4003), .ZN(n2490) );
  NOR2_X2 U2813 ( .A1(n2528), .A2(n4242), .ZN(n4274) );
  INV_X4 U2814 ( .A(n2410), .ZN(n1041) );
  OR2_X2 U2815 ( .A1(n4401), .A2(n4516), .ZN(n2719) );
  INV_X2 U2817 ( .A(n4257), .ZN(n4227) );
  NOR2_X2 U2818 ( .A1(n5269), .A2(n5268), .ZN(n5273) );
  INV_X1 U2819 ( .A(n4162), .ZN(n4192) );
  INV_X2 U2821 ( .A(n4139), .ZN(n4145) );
  NAND2_X1 U2822 ( .A1(n4140), .A2(n4141), .ZN(n4144) );
  INV_X2 U2825 ( .A(n5949), .ZN(n5950) );
  NAND2_X2 U2828 ( .A1(n3784), .A2(n3783), .ZN(n3814) );
  NAND2_X1 U2829 ( .A1(n6047), .A2(n6038), .ZN(n6036) );
  INV_X4 U2830 ( .A(n3571), .ZN(n1043) );
  NOR2_X1 U2832 ( .A1(n6047), .A2(n6046), .ZN(n6102) );
  INV_X4 U2834 ( .A(n3885), .ZN(n1046) );
  INV_X2 U2836 ( .A(n4796), .ZN(n1464) );
  INV_X4 U2837 ( .A(n4451), .ZN(n1047) );
  AOI22_X1 U2839 ( .A1(n3351), .A2(n5951), .B1(n5471), .B2(n5526), .ZN(n1618)
         );
  NAND2_X1 U2840 ( .A1(b[0]), .A2(n6215), .ZN(n4126) );
  NAND2_X1 U2841 ( .A1(n6045), .A2(n6044), .ZN(n6046) );
  INV_X4 U2843 ( .A(n5283), .ZN(n1048) );
  INV_X2 U2845 ( .A(n2027), .ZN(n2028) );
  INV_X2 U2846 ( .A(n4032), .ZN(n1049) );
  INV_X4 U2847 ( .A(n3890), .ZN(n1050) );
  INV_X4 U2850 ( .A(n3802), .ZN(n1051) );
  INV_X2 U2851 ( .A(n5228), .ZN(n5225) );
  INV_X4 U2852 ( .A(n4099), .ZN(n1052) );
  INV_X2 U2853 ( .A(n4121), .ZN(n4123) );
  AOI21_X1 U2854 ( .B1(n6043), .B2(b[23]), .A(n6042), .ZN(n6044) );
  INV_X2 U2859 ( .A(n4245), .ZN(n4246) );
  INV_X2 U2861 ( .A(n4237), .ZN(n4241) );
  NAND2_X2 U2862 ( .A1(n2197), .A2(n2196), .ZN(n3888) );
  NOR3_X2 U2863 ( .A1(n2462), .A2(n6160), .A3(n3756), .ZN(n2463) );
  INV_X4 U2864 ( .A(n4936), .ZN(n1055) );
  AND2_X2 U2865 ( .A1(n5106), .A2(b[13]), .ZN(n3761) );
  INV_X1 U2866 ( .A(n6041), .ZN(n6042) );
  INV_X2 U2867 ( .A(n4378), .ZN(n3971) );
  INV_X2 U2869 ( .A(n4189), .ZN(n1058) );
  NAND2_X2 U2871 ( .A1(n441), .A2(b[1]), .ZN(n1686) );
  INV_X2 U2872 ( .A(n4133), .ZN(n6096) );
  NAND2_X1 U2873 ( .A1(n6033), .A2(b[21]), .ZN(n6041) );
  INV_X2 U2874 ( .A(n4697), .ZN(n4698) );
  INV_X8 U2875 ( .A(n3484), .ZN(n1059) );
  NOR2_X1 U2876 ( .A1(n4783), .A2(n4784), .ZN(n2885) );
  INV_X2 U2878 ( .A(n5957), .ZN(n6033) );
  NAND2_X2 U2879 ( .A1(n5957), .A2(n5951), .ZN(n6038) );
  OR2_X2 U2883 ( .A1(n5952), .A2(b[6]), .ZN(n2734) );
  INV_X2 U2884 ( .A(n4846), .ZN(n1061) );
  AND2_X2 U2886 ( .A1(n2045), .A2(a[17]), .ZN(n5422) );
  INV_X2 U2887 ( .A(n5531), .ZN(n5516) );
  NOR2_X1 U2888 ( .A1(n2032), .A2(a[17]), .ZN(n5409) );
  XNOR2_X1 U2890 ( .A(a[13]), .B(b[3]), .ZN(n2716) );
  OR2_X2 U2892 ( .A1(a[19]), .A2(a[20]), .ZN(n3762) );
  INV_X4 U2893 ( .A(n4834), .ZN(n1062) );
  XNOR2_X1 U2894 ( .A(a[17]), .B(b[6]), .ZN(n4417) );
  XOR2_X2 U2895 ( .A(a[7]), .B(b[15]), .Z(n4321) );
  OAI21_X1 U2896 ( .B1(b[15]), .B2(b[14]), .A(a[23]), .ZN(n5469) );
  XNOR2_X1 U2897 ( .A(a[11]), .B(b[5]), .ZN(n3854) );
  XOR2_X2 U2899 ( .A(b[7]), .B(a[21]), .Z(n4742) );
  XNOR2_X1 U2901 ( .A(a[9]), .B(b[5]), .ZN(n3795) );
  XOR2_X2 U2902 ( .A(a[1]), .B(b[13]), .Z(n3809) );
  XNOR2_X1 U2907 ( .A(b[15]), .B(b[14]), .ZN(n5498) );
  NAND2_X2 U2911 ( .A1(a[23]), .A2(b[14]), .ZN(n5450) );
  XNOR2_X1 U2913 ( .A(a[17]), .B(b[5]), .ZN(n4355) );
  XOR2_X2 U2915 ( .A(a[15]), .B(b[17]), .Z(n4922) );
  XNOR2_X1 U2916 ( .A(a[7]), .B(b[20]), .ZN(n4693) );
  INV_X1 U2918 ( .A(b[20]), .ZN(n3372) );
  INV_X2 U2919 ( .A(b[7]), .ZN(n2143) );
  NAND2_X1 U2920 ( .A1(b[17]), .A2(b[16]), .ZN(n5397) );
  XNOR2_X1 U2921 ( .A(b[7]), .B(a[9]), .ZN(n3849) );
  XOR2_X2 U2926 ( .A(a[15]), .B(b[14]), .Z(n4847) );
  XNOR2_X1 U2928 ( .A(b[12]), .B(a[19]), .ZN(n4896) );
  OAI21_X1 U2929 ( .B1(b[18]), .B2(b[19]), .A(a[23]), .ZN(n5904) );
  XOR2_X2 U2930 ( .A(a[17]), .B(b[19]), .Z(n5168) );
  INV_X4 U2932 ( .A(b[17]), .ZN(n3217) );
  NAND2_X2 U2933 ( .A1(n4242), .A2(n2528), .ZN(n4276) );
  NAND2_X2 U2935 ( .A1(n1065), .A2(n1256), .ZN(n2193) );
  NOR2_X2 U2936 ( .A1(n3503), .A2(n531), .ZN(n1065) );
  INV_X4 U2937 ( .A(n5086), .ZN(n5089) );
  BUF_X4 U2939 ( .A(n4886), .Z(n1207) );
  NAND2_X1 U2940 ( .A1(n4920), .A2(n4921), .ZN(n2751) );
  INV_X4 U2941 ( .A(n2029), .ZN(n3627) );
  NAND2_X2 U2943 ( .A1(n3302), .A2(n3303), .ZN(n4472) );
  BUF_X4 U2946 ( .A(n1089), .Z(n1067) );
  NAND2_X2 U2947 ( .A1(n1089), .A2(n4969), .ZN(n5809) );
  NAND2_X2 U2949 ( .A1(n1696), .A2(n4668), .ZN(n1068) );
  NAND2_X2 U2950 ( .A1(n1072), .A2(n1071), .ZN(n1696) );
  NAND2_X2 U2951 ( .A1(n1338), .A2(n1030), .ZN(n1072) );
  NAND3_X2 U2952 ( .A1(n1417), .A2(n1074), .A3(n1073), .ZN(n2787) );
  NAND2_X1 U2953 ( .A1(n1653), .A2(n1844), .ZN(n1074) );
  NAND2_X2 U2954 ( .A1(n1848), .A2(n2787), .ZN(n1084) );
  INV_X4 U2955 ( .A(n4616), .ZN(n4619) );
  NAND2_X4 U2956 ( .A1(b[0]), .A2(a[23]), .ZN(n4616) );
  XNOR2_X2 U2957 ( .A(n4617), .B(n4619), .ZN(n2459) );
  OAI21_X2 U2958 ( .B1(n1075), .B2(a[0]), .A(a[1]), .ZN(n4617) );
  NAND4_X1 U2959 ( .A1(n5809), .A2(n3672), .A3(n6093), .A4(n6092), .ZN(n3770)
         );
  NAND2_X2 U2960 ( .A1(n1663), .A2(n1664), .ZN(n4969) );
  NAND3_X1 U2961 ( .A1(n1848), .A2(n2787), .A3(n2391), .ZN(n1080) );
  NAND2_X2 U2962 ( .A1(n1084), .A2(n1082), .ZN(n1081) );
  BUF_X4 U2963 ( .A(n3126), .Z(n1085) );
  NOR2_X1 U2964 ( .A1(n5804), .A2(n3126), .ZN(n4986) );
  NAND2_X2 U2965 ( .A1(n1088), .A2(n1086), .ZN(n1522) );
  XNOR2_X2 U2967 ( .A(n1087), .B(n459), .ZN(n4881) );
  XNOR2_X2 U2970 ( .A(n1336), .B(n1950), .ZN(n3468) );
  NAND3_X2 U2971 ( .A1(n1249), .A2(n1254), .A3(n1335), .ZN(n2571) );
  NAND3_X2 U2974 ( .A1(n4657), .A2(n2215), .A3(n3648), .ZN(n2548) );
  NOR2_X2 U2977 ( .A1(n5839), .A2(n4986), .ZN(n4987) );
  INV_X4 U2978 ( .A(n1235), .ZN(n1857) );
  NAND2_X2 U2979 ( .A1(n1090), .A2(n2751), .ZN(n1619) );
  NAND2_X2 U2980 ( .A1(n2753), .A2(n2752), .ZN(n1090) );
  NAND2_X2 U2981 ( .A1(n1092), .A2(n1091), .ZN(n1164) );
  NAND2_X2 U2982 ( .A1(n4483), .A2(b[7]), .ZN(n1092) );
  NAND2_X2 U2983 ( .A1(n3596), .A2(n3155), .ZN(n3316) );
  NAND2_X2 U2984 ( .A1(n1024), .A2(n1025), .ZN(n1301) );
  NAND2_X2 U2985 ( .A1(n6622), .A2(n4737), .ZN(n2022) );
  NAND2_X2 U2986 ( .A1(n2024), .A2(n6351), .ZN(n4739) );
  AOI21_X2 U2987 ( .B1(n2326), .B2(n2723), .A(n1208), .ZN(n4002) );
  NAND2_X4 U2988 ( .A1(n1854), .A2(n1094), .ZN(n1119) );
  NAND3_X2 U2989 ( .A1(n1853), .A2(n1235), .A3(n4685), .ZN(n1094) );
  NAND2_X2 U2994 ( .A1(n2530), .A2(n4487), .ZN(n2120) );
  AOI21_X2 U2995 ( .B1(n320), .B2(n4044), .A(n3322), .ZN(n4465) );
  INV_X4 U2997 ( .A(n1799), .ZN(n1803) );
  INV_X2 U2998 ( .A(n3350), .ZN(n1744) );
  NOR2_X4 U2999 ( .A1(n3704), .A2(n4500), .ZN(n2487) );
  INV_X2 U3002 ( .A(n2612), .ZN(n2611) );
  NAND2_X2 U3003 ( .A1(n4578), .A2(n4577), .ZN(n2612) );
  BUF_X4 U3005 ( .A(n4285), .Z(n1097) );
  INV_X4 U3007 ( .A(n2310), .ZN(n3743) );
  NOR2_X2 U3009 ( .A1(n1655), .A2(n1485), .ZN(n3376) );
  BUF_X4 U3010 ( .A(n5919), .Z(n1099) );
  NAND2_X2 U3011 ( .A1(n3173), .A2(n3174), .ZN(n2299) );
  NAND2_X2 U3012 ( .A1(n2111), .A2(n2110), .ZN(n3173) );
  INV_X4 U3014 ( .A(n3674), .ZN(n4526) );
  NOR2_X4 U3015 ( .A1(n5570), .A2(n5571), .ZN(n5999) );
  NAND2_X2 U3016 ( .A1(n1102), .A2(n1101), .ZN(n4433) );
  NAND2_X2 U3017 ( .A1(n4774), .A2(b[8]), .ZN(n1101) );
  AOI22_X2 U3018 ( .A1(n5277), .A2(n435), .B1(b[12]), .B2(n5900), .ZN(n5192)
         );
  INV_X4 U3021 ( .A(n1005), .ZN(n2491) );
  INV_X4 U3023 ( .A(n3704), .ZN(n2103) );
  NOR2_X4 U3025 ( .A1(n3773), .A2(n635), .ZN(n4238) );
  AOI22_X2 U3026 ( .A1(n3701), .A2(n1106), .B1(n2565), .B2(n1626), .ZN(n2564)
         );
  NOR2_X2 U3027 ( .A1(n1626), .A2(n4084), .ZN(n1106) );
  OAI21_X2 U3028 ( .B1(n2596), .B2(n2595), .A(n4789), .ZN(n4840) );
  NOR3_X4 U3029 ( .A1(n4156), .A2(n4155), .A3(n4154), .ZN(n3722) );
  NAND2_X2 U3031 ( .A1(n2896), .A2(n2897), .ZN(n1835) );
  INV_X4 U3032 ( .A(n1281), .ZN(n3202) );
  NAND3_X2 U3033 ( .A1(n4751), .A2(n4846), .A3(n5190), .ZN(n3280) );
  NOR3_X4 U3035 ( .A1(n3684), .A2(a[7]), .A3(a[8]), .ZN(n4795) );
  BUF_X4 U3036 ( .A(n6326), .Z(n1107) );
  NAND2_X2 U3037 ( .A1(n1109), .A2(n1108), .ZN(n4951) );
  NAND2_X2 U3038 ( .A1(n2382), .A2(b[14]), .ZN(n1108) );
  NAND2_X2 U3039 ( .A1(n2510), .A2(n5293), .ZN(n1109) );
  INV_X4 U3041 ( .A(n2226), .ZN(n2708) );
  NOR2_X2 U3042 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  INV_X4 U3043 ( .A(n4902), .ZN(n2628) );
  INV_X4 U3045 ( .A(n3561), .ZN(n2081) );
  NOR2_X4 U3047 ( .A1(n3909), .A2(a[17]), .ZN(n5423) );
  NAND2_X2 U3048 ( .A1(n5039), .A2(n3074), .ZN(n1112) );
  NAND2_X2 U3049 ( .A1(n1114), .A2(n1113), .ZN(n2058) );
  NAND2_X2 U3050 ( .A1(b[10]), .A2(n4483), .ZN(n1114) );
  INV_X8 U3054 ( .A(a[23]), .ZN(n5952) );
  OAI21_X2 U3055 ( .B1(n1116), .B2(n2377), .A(n2376), .ZN(n4232) );
  NAND2_X2 U3057 ( .A1(n5694), .A2(n5689), .ZN(n1118) );
  NAND2_X2 U3058 ( .A1(n1118), .A2(n1117), .ZN(n4195) );
  OAI21_X2 U3059 ( .B1(n4671), .B2(n1119), .A(n1851), .ZN(n2231) );
  XNOR2_X2 U3060 ( .A(n1119), .B(n3755), .ZN(n1239) );
  NAND2_X4 U3064 ( .A1(a[4]), .A2(a[3]), .ZN(n1121) );
  XNOR2_X2 U3068 ( .A(n3034), .B(n4261), .ZN(n1125) );
  XNOR2_X2 U3069 ( .A(n1126), .B(n4227), .ZN(n4261) );
  NAND3_X2 U3072 ( .A1(n4215), .A2(n2186), .A3(n2185), .ZN(n4308) );
  INV_X4 U3074 ( .A(n3617), .ZN(n1127) );
  AOI21_X2 U3075 ( .B1(n1130), .B2(n1129), .A(n1128), .ZN(n4152) );
  INV_X2 U3076 ( .A(n4098), .ZN(n1130) );
  NAND2_X2 U3077 ( .A1(n1789), .A2(n1131), .ZN(n1786) );
  XNOR2_X2 U3079 ( .A(n1789), .B(n1131), .ZN(n1222) );
  NAND2_X4 U3080 ( .A1(n1303), .A2(n1304), .ZN(n1131) );
  INV_X4 U3081 ( .A(n1132), .ZN(n3470) );
  NAND2_X4 U3082 ( .A1(n2035), .A2(n2036), .ZN(n1132) );
  NOR2_X2 U3083 ( .A1(n5671), .A2(n4206), .ZN(n1133) );
  NAND2_X2 U3084 ( .A1(n4203), .A2(n4202), .ZN(n5671) );
  NOR2_X2 U3085 ( .A1(n1135), .A2(n5676), .ZN(n1134) );
  AOI21_X2 U3086 ( .B1(n4203), .B2(n4200), .A(n5675), .ZN(n1135) );
  AOI21_X2 U3087 ( .B1(n545), .B2(n4196), .A(n1770), .ZN(n5675) );
  INV_X4 U3088 ( .A(n4228), .ZN(n4187) );
  AOI21_X2 U3089 ( .B1(n6558), .B2(n4186), .A(n4185), .ZN(n4228) );
  NAND2_X2 U3090 ( .A1(n4231), .A2(n2508), .ZN(n1138) );
  NAND2_X2 U3091 ( .A1(n2604), .A2(b[1]), .ZN(n1139) );
  NAND2_X2 U3093 ( .A1(n1143), .A2(n4714), .ZN(\d[26]_BAR ) );
  INV_X2 U3094 ( .A(n1144), .ZN(n1143) );
  NAND2_X2 U3095 ( .A1(n600), .A2(n6013), .ZN(n6020) );
  NAND2_X2 U3098 ( .A1(n1147), .A2(b[18]), .ZN(n2592) );
  NAND2_X2 U3099 ( .A1(n1147), .A2(b[1]), .ZN(n3592) );
  NOR2_X1 U3102 ( .A1(n711), .A2(n4475), .ZN(n1153) );
  NAND2_X2 U3104 ( .A1(n4472), .A2(n2865), .ZN(n2118) );
  NAND2_X1 U3105 ( .A1(n3569), .A2(n4374), .ZN(n1158) );
  NAND2_X2 U3106 ( .A1(n2088), .A2(n2907), .ZN(n1159) );
  INV_X2 U3107 ( .A(n2937), .ZN(n3297) );
  NAND2_X2 U3108 ( .A1(n964), .A2(n4554), .ZN(n1160) );
  OAI21_X2 U3109 ( .B1(n964), .B2(n4554), .A(n4555), .ZN(n1161) );
  NAND2_X2 U3111 ( .A1(n4761), .A2(n4760), .ZN(n1578) );
  NAND3_X2 U3113 ( .A1(n1165), .A2(n1580), .A3(n1167), .ZN(n4761) );
  NAND2_X2 U3114 ( .A1(n962), .A2(n1166), .ZN(n1580) );
  NAND2_X2 U3115 ( .A1(n4696), .A2(n4933), .ZN(n1165) );
  INV_X8 U3116 ( .A(n3395), .ZN(n4933) );
  INV_X2 U3117 ( .A(n4045), .ZN(n1166) );
  AOI22_X2 U3119 ( .A1(n4695), .A2(n4998), .B1(a[9]), .B2(b[18]), .ZN(n4696)
         );
  INV_X2 U3120 ( .A(n1168), .ZN(n2674) );
  NOR2_X2 U3121 ( .A1(n3545), .A2(n4763), .ZN(n1168) );
  NAND2_X2 U3122 ( .A1(n1170), .A2(n1169), .ZN(n4858) );
  NAND2_X2 U3124 ( .A1(n1172), .A2(n1171), .ZN(n1170) );
  NAND2_X2 U3126 ( .A1(n2392), .A2(n4840), .ZN(n1172) );
  NAND2_X2 U3127 ( .A1(n1726), .A2(n1725), .ZN(n2392) );
  INV_X2 U3128 ( .A(n3986), .ZN(n1174) );
  NAND2_X2 U3129 ( .A1(n2208), .A2(n6359), .ZN(n1175) );
  XNOR2_X2 U3130 ( .A(n2209), .B(n2210), .ZN(n3984) );
  NAND2_X2 U3131 ( .A1(n1174), .A2(n1173), .ZN(n2669) );
  INV_X2 U3134 ( .A(n1178), .ZN(n5465) );
  NAND2_X2 U3135 ( .A1(n5503), .A2(n1179), .ZN(n1178) );
  NAND2_X2 U3136 ( .A1(n5448), .A2(n5460), .ZN(n5503) );
  AOI21_X2 U3137 ( .B1(n5447), .B2(n5496), .A(n5495), .ZN(n5460) );
  NAND2_X2 U3138 ( .A1(n3486), .A2(n3485), .ZN(n5448) );
  NAND2_X2 U3140 ( .A1(n1181), .A2(n1182), .ZN(n3480) );
  NAND3_X1 U3141 ( .A1(n1182), .A2(n4918), .A3(n1181), .ZN(n3077) );
  NAND2_X2 U3143 ( .A1(n2847), .A2(n1954), .ZN(n1182) );
  BUF_X4 U3144 ( .A(n3480), .Z(n1183) );
  INV_X1 U3145 ( .A(n487), .ZN(n5035) );
  NAND2_X1 U3146 ( .A1(n5031), .A2(n487), .ZN(n5033) );
  NAND2_X2 U3148 ( .A1(n3326), .A2(n3572), .ZN(n1185) );
  INV_X4 U3149 ( .A(n1186), .ZN(n2281) );
  NAND2_X2 U3150 ( .A1(n2995), .A2(n1717), .ZN(n1186) );
  NAND3_X2 U3151 ( .A1(n2474), .A2(n1186), .A3(n3714), .ZN(n3712) );
  INV_X2 U3152 ( .A(n2802), .ZN(n4902) );
  NAND2_X2 U3154 ( .A1(n2028), .A2(n2026), .ZN(n4731) );
  NAND2_X2 U3155 ( .A1(n4730), .A2(n4732), .ZN(n1689) );
  INV_X2 U3156 ( .A(n4728), .ZN(n4729) );
  INV_X2 U3157 ( .A(n1187), .ZN(n1609) );
  NAND2_X2 U3158 ( .A1(n1188), .A2(n1187), .ZN(n5573) );
  NAND2_X2 U3159 ( .A1(n1612), .A2(n1608), .ZN(n1187) );
  INV_X2 U3160 ( .A(n1610), .ZN(n1188) );
  INV_X2 U3161 ( .A(n5425), .ZN(n1190) );
  OAI21_X2 U3162 ( .B1(n5424), .B2(n5425), .A(n1189), .ZN(n3488) );
  INV_X1 U3163 ( .A(n3488), .ZN(n5436) );
  AOI21_X2 U3164 ( .B1(n5437), .B2(n3488), .A(n5438), .ZN(n3487) );
  NOR3_X2 U3165 ( .A1(n3440), .A2(n5426), .A3(n3441), .ZN(n5438) );
  NAND2_X2 U3166 ( .A1(n1196), .A2(n1195), .ZN(n1192) );
  BUF_X4 U3167 ( .A(n4768), .Z(n1193) );
  NAND2_X2 U3168 ( .A1(n5454), .A2(b[14]), .ZN(n1196) );
  OAI21_X2 U3169 ( .B1(n1198), .B2(n2013), .A(n4562), .ZN(n1197) );
  INV_X2 U3170 ( .A(n1199), .ZN(n1198) );
  NAND2_X2 U3173 ( .A1(n442), .A2(n443), .ZN(n2178) );
  NAND2_X2 U3176 ( .A1(n1203), .A2(n3752), .ZN(n2979) );
  NOR2_X2 U3177 ( .A1(n1203), .A2(n3752), .ZN(n2980) );
  INV_X4 U3178 ( .A(n2825), .ZN(n1203) );
  AOI21_X2 U3179 ( .B1(n2074), .B2(n1205), .A(n1204), .ZN(n5171) );
  XNOR2_X2 U3183 ( .A(n4003), .B(n4002), .ZN(n2545) );
  OAI21_X2 U3185 ( .B1(n3795), .B2(n3617), .A(n1209), .ZN(n4003) );
  NAND2_X2 U3186 ( .A1(n1211), .A2(n1210), .ZN(n1209) );
  NAND2_X2 U3187 ( .A1(n4810), .A2(b[4]), .ZN(n1211) );
  NOR2_X2 U3188 ( .A1(n4694), .A2(n1212), .ZN(n2737) );
  INV_X2 U3189 ( .A(b[17]), .ZN(n1212) );
  NAND2_X2 U3190 ( .A1(n1213), .A2(a[7]), .ZN(n4694) );
  INV_X2 U3191 ( .A(a[9]), .ZN(n1213) );
  NAND2_X2 U3195 ( .A1(n1217), .A2(n4852), .ZN(n4864) );
  AOI22_X2 U3196 ( .A1(n1218), .A2(n4844), .B1(n5010), .B2(n4843), .ZN(n4852)
         );
  INV_X2 U3197 ( .A(n1219), .ZN(n1217) );
  INV_X2 U3198 ( .A(n5899), .ZN(n5948) );
  INV_X2 U3201 ( .A(n4860), .ZN(n1221) );
  AOI21_X2 U3202 ( .B1(n4907), .B2(n4908), .A(n4916), .ZN(n3680) );
  NOR2_X4 U3203 ( .A1(n994), .A2(n2311), .ZN(n4916) );
  NAND3_X2 U3204 ( .A1(n1956), .A2(n2349), .A3(n2348), .ZN(n1223) );
  INV_X4 U3205 ( .A(n1226), .ZN(n2351) );
  NAND2_X2 U3206 ( .A1(n2492), .A2(n3411), .ZN(n1226) );
  AOI22_X2 U3207 ( .A1(n1227), .A2(n957), .B1(n2316), .B2(n2978), .ZN(n3411)
         );
  INV_X2 U3208 ( .A(n2312), .ZN(n1227) );
  NAND2_X2 U3209 ( .A1(n1228), .A2(n4833), .ZN(n2492) );
  OAI21_X2 U3212 ( .B1(n1231), .B2(n4838), .A(n1229), .ZN(n4914) );
  NAND2_X2 U3213 ( .A1(n2351), .A2(n2350), .ZN(n1229) );
  NOR2_X2 U3214 ( .A1(n2350), .A2(n2351), .ZN(n1231) );
  NAND2_X2 U3218 ( .A1(n3752), .A2(n2825), .ZN(n1235) );
  NAND2_X4 U3219 ( .A1(n1236), .A2(n2001), .ZN(n2384) );
  NAND2_X2 U3220 ( .A1(n3283), .A2(n6449), .ZN(n1236) );
  NAND2_X2 U3222 ( .A1(n2802), .A2(n3250), .ZN(n1555) );
  NOR2_X1 U3223 ( .A1(n2244), .A2(n3367), .ZN(n1767) );
  NOR2_X1 U3224 ( .A1(n2244), .A2(n3835), .ZN(n3837) );
  NAND2_X1 U3225 ( .A1(n2244), .A2(b[15]), .ZN(n3328) );
  NAND2_X1 U3226 ( .A1(n2244), .A2(b[13]), .ZN(n4336) );
  NAND2_X1 U3227 ( .A1(n2244), .A2(b[14]), .ZN(n2413) );
  NAND2_X1 U3228 ( .A1(n2244), .A2(b[16]), .ZN(n2145) );
  AOI22_X1 U3231 ( .A1(n3342), .A2(n1847), .B1(n2244), .B2(b[8]), .ZN(n3228)
         );
  AOI22_X2 U3232 ( .A1(n2678), .A2(n2679), .B1(n3150), .B2(n4803), .ZN(n3313)
         );
  XNOR2_X2 U3233 ( .A(n1440), .B(n4883), .ZN(n1242) );
  NOR2_X4 U3234 ( .A1(n2529), .A2(n4583), .ZN(n2681) );
  NAND2_X2 U3235 ( .A1(n1244), .A2(n1017), .ZN(n1243) );
  NAND2_X1 U3236 ( .A1(n4473), .A2(n1754), .ZN(n1244) );
  NAND2_X2 U3239 ( .A1(n1247), .A2(n2601), .ZN(n1246) );
  NOR3_X4 U3240 ( .A1(n1248), .A2(a[1]), .A3(a[2]), .ZN(n4543) );
  INV_X8 U3241 ( .A(a[3]), .ZN(n1248) );
  NAND2_X2 U3242 ( .A1(n2193), .A2(n2192), .ZN(n1795) );
  NAND3_X2 U3243 ( .A1(n1960), .A2(n2399), .A3(n1062), .ZN(n1252) );
  INV_X2 U3244 ( .A(n4835), .ZN(n1255) );
  NAND2_X4 U3246 ( .A1(n6615), .A2(a[11]), .ZN(n4886) );
  NOR2_X4 U3247 ( .A1(a[9]), .A2(a[10]), .ZN(n3991) );
  NAND3_X2 U3249 ( .A1(n3947), .A2(n3626), .A3(n3940), .ZN(n1257) );
  NAND2_X2 U3250 ( .A1(n3297), .A2(n2939), .ZN(n1258) );
  INV_X4 U3256 ( .A(n2898), .ZN(n2775) );
  NAND2_X2 U3257 ( .A1(n647), .A2(n1263), .ZN(n2898) );
  XNOR2_X2 U3259 ( .A(n3232), .B(n6193), .ZN(n1265) );
  NAND2_X4 U3260 ( .A1(n1287), .A2(n2713), .ZN(n3251) );
  NAND2_X2 U3261 ( .A1(n3251), .A2(n3386), .ZN(n2315) );
  NOR2_X2 U3264 ( .A1(n1271), .A2(n1045), .ZN(n1270) );
  INV_X2 U3265 ( .A(n5052), .ZN(n1271) );
  OAI21_X2 U3266 ( .B1(n5004), .B2(n5005), .A(n1625), .ZN(n1272) );
  NOR2_X2 U3269 ( .A1(n3704), .A2(n5003), .ZN(n5004) );
  NAND2_X2 U3270 ( .A1(n5054), .A2(n5053), .ZN(n1273) );
  OAI21_X2 U3273 ( .B1(n4038), .B2(n4037), .A(n3594), .ZN(n1275) );
  XNOR2_X2 U3275 ( .A(n4612), .B(n4562), .ZN(n2177) );
  NAND2_X2 U3276 ( .A1(n4564), .A2(n4563), .ZN(n1279) );
  AOI22_X2 U3277 ( .A1(n969), .A2(n781), .B1(n780), .B2(n1003), .ZN(n1822) );
  OAI21_X2 U3279 ( .B1(n4076), .B2(n4077), .A(n4075), .ZN(n3615) );
  NAND2_X2 U3280 ( .A1(n3108), .A2(n759), .ZN(n1377) );
  NAND3_X2 U3281 ( .A1(n6516), .A2(n1283), .A3(n3628), .ZN(n3108) );
  NAND2_X2 U3282 ( .A1(n3106), .A2(n2029), .ZN(n3629) );
  AOI22_X2 U3284 ( .A1(n3644), .A2(n3643), .B1(n3763), .B2(n1287), .ZN(n3268)
         );
  INV_X8 U3285 ( .A(n4776), .ZN(n1287) );
  AOI22_X2 U3286 ( .A1(n4397), .A2(n3328), .B1(n1287), .B2(n4398), .ZN(n4509)
         );
  NAND2_X2 U3288 ( .A1(n2718), .A2(n1287), .ZN(n3227) );
  NAND2_X2 U3289 ( .A1(n4689), .A2(n1287), .ZN(n4236) );
  AOI22_X2 U3291 ( .A1(n2145), .A2(n2146), .B1(n4482), .B2(n1287), .ZN(n4567)
         );
  AOI22_X2 U3292 ( .A1(n4336), .A2(n4335), .B1(n4334), .B2(n1287), .ZN(n4382)
         );
  BUF_X4 U3293 ( .A(n1547), .Z(n1288) );
  NAND2_X2 U3294 ( .A1(n1289), .A2(n3981), .ZN(n2298) );
  NAND2_X1 U3295 ( .A1(n3983), .A2(n1289), .ZN(n1401) );
  INV_X4 U3298 ( .A(n1291), .ZN(n1290) );
  NOR2_X2 U3299 ( .A1(n3911), .A2(n1056), .ZN(n1291) );
  NAND2_X2 U3300 ( .A1(n1293), .A2(n2308), .ZN(n1292) );
  NOR2_X2 U3306 ( .A1(n3189), .A2(n3188), .ZN(n1302) );
  NAND2_X2 U3307 ( .A1(n1301), .A2(n1300), .ZN(n3189) );
  INV_X2 U3308 ( .A(n1302), .ZN(n2080) );
  NAND2_X2 U3309 ( .A1(n1577), .A2(n1576), .ZN(n1303) );
  NAND2_X2 U3310 ( .A1(n1578), .A2(n4762), .ZN(n1304) );
  XNOR2_X2 U3311 ( .A(a[17]), .B(b[10]), .ZN(n4709) );
  NAND2_X2 U3312 ( .A1(n2109), .A2(n3190), .ZN(n3174) );
  NAND3_X2 U3313 ( .A1(n1953), .A2(n584), .A3(n2003), .ZN(n1305) );
  NAND2_X2 U3314 ( .A1(n4879), .A2(n4878), .ZN(n4880) );
  NAND2_X2 U3315 ( .A1(n6327), .A2(n3113), .ZN(n4879) );
  INV_X4 U3318 ( .A(n2171), .ZN(n2436) );
  BUF_X4 U3319 ( .A(n3461), .Z(n1307) );
  BUF_X4 U3320 ( .A(n1847), .Z(n1308) );
  BUF_X4 U3321 ( .A(n5681), .Z(n1309) );
  NAND4_X1 U3323 ( .A1(n2118), .A2(n2120), .A3(n6149), .A4(n2119), .ZN(n2168)
         );
  NAND2_X2 U3324 ( .A1(n1311), .A2(n2665), .ZN(n2059) );
  NAND2_X2 U3325 ( .A1(n1313), .A2(n1312), .ZN(n1311) );
  INV_X2 U3326 ( .A(n5565), .ZN(n1312) );
  INV_X2 U3327 ( .A(n2861), .ZN(n1313) );
  BUF_X4 U3328 ( .A(n6005), .Z(n1314) );
  BUF_X4 U3329 ( .A(n5676), .Z(n1315) );
  NOR2_X4 U3330 ( .A1(n3820), .A2(n3819), .ZN(n3858) );
  NAND2_X2 U3331 ( .A1(n1316), .A2(n2664), .ZN(n3518) );
  NAND2_X2 U3332 ( .A1(n2662), .A2(n2663), .ZN(n1316) );
  NAND2_X2 U3333 ( .A1(n1750), .A2(n1317), .ZN(n1751) );
  NAND2_X2 U3334 ( .A1(n2061), .A2(n2060), .ZN(n2064) );
  NAND3_X2 U3335 ( .A1(n3039), .A2(n4250), .A3(n3040), .ZN(n2185) );
  NAND2_X2 U3336 ( .A1(n4672), .A2(n3268), .ZN(n1938) );
  NAND2_X2 U3337 ( .A1(n1048), .A2(n1037), .ZN(n2661) );
  NAND2_X2 U3338 ( .A1(n4934), .A2(n4933), .ZN(n2586) );
  OAI21_X2 U3339 ( .B1(n5027), .B2(n5028), .A(n1035), .ZN(n2477) );
  AOI21_X2 U3341 ( .B1(n1425), .B2(n5155), .A(n5154), .ZN(n5212) );
  AOI22_X2 U3342 ( .A1(n258), .A2(n2655), .B1(n5089), .B2(n5088), .ZN(n5155)
         );
  OAI21_X2 U3343 ( .B1(n6506), .B2(n3149), .A(n3220), .ZN(n1850) );
  BUF_X4 U3344 ( .A(n2037), .Z(n1318) );
  NAND2_X2 U3346 ( .A1(n3012), .A2(n5621), .ZN(n5160) );
  NAND2_X2 U3347 ( .A1(n1374), .A2(n5383), .ZN(n5621) );
  NOR2_X4 U3348 ( .A1(n2774), .A2(n3200), .ZN(n2931) );
  AOI21_X2 U3349 ( .B1(n4285), .B2(n3582), .A(n4284), .ZN(n2438) );
  BUF_X4 U3354 ( .A(n4299), .Z(n1320) );
  NAND2_X2 U3355 ( .A1(n5817), .A2(n2087), .ZN(n3520) );
  NAND2_X2 U3356 ( .A1(n1600), .A2(n1601), .ZN(n5817) );
  INV_X2 U3359 ( .A(n1923), .ZN(n1321) );
  NOR2_X4 U3361 ( .A1(n3699), .A2(n4400), .ZN(n4516) );
  NAND2_X2 U3362 ( .A1(n3132), .A2(n1322), .ZN(n4510) );
  OAI21_X2 U3364 ( .B1(n4877), .B2(n46), .A(n4875), .ZN(n4892) );
  NAND2_X2 U3367 ( .A1(n1325), .A2(n1323), .ZN(n3805) );
  NAND2_X2 U3368 ( .A1(n1308), .A2(n1324), .ZN(n1323) );
  NAND2_X2 U3369 ( .A1(n6203), .A2(b[6]), .ZN(n1325) );
  AOI21_X2 U3370 ( .B1(n1986), .B2(n4912), .A(n1940), .ZN(n3608) );
  NAND2_X2 U3371 ( .A1(n2080), .A2(n2079), .ZN(n4910) );
  NOR2_X2 U3372 ( .A1(n5707), .A2(n5704), .ZN(n2364) );
  NAND2_X2 U3374 ( .A1(n1326), .A2(n3261), .ZN(n1501) );
  NOR2_X2 U3376 ( .A1(n2822), .A2(n3724), .ZN(n1327) );
  NOR2_X2 U3377 ( .A1(n1328), .A2(n3585), .ZN(n2008) );
  NAND2_X2 U3378 ( .A1(n2895), .A2(n2948), .ZN(n1328) );
  NOR2_X4 U3379 ( .A1(n6589), .A2(n4828), .ZN(n1591) );
  OAI21_X2 U3380 ( .B1(n1331), .B2(n3066), .A(n1330), .ZN(n1531) );
  INV_X8 U3383 ( .A(n6459), .ZN(n3704) );
  NAND3_X2 U3384 ( .A1(n1635), .A2(n1636), .A3(n5033), .ZN(n1634) );
  NAND2_X2 U3385 ( .A1(n2320), .A2(n3682), .ZN(n3681) );
  NOR2_X2 U3386 ( .A1(n6511), .A2(n4964), .ZN(n3379) );
  INV_X4 U3390 ( .A(n3408), .ZN(n2144) );
  NAND2_X2 U3391 ( .A1(n1334), .A2(n1018), .ZN(n2040) );
  NAND2_X2 U3393 ( .A1(n4833), .A2(n3412), .ZN(n1335) );
  NOR2_X4 U3394 ( .A1(n3345), .A2(n2533), .ZN(n4020) );
  NAND2_X2 U3396 ( .A1(n699), .A2(n4942), .ZN(n3576) );
  INV_X4 U3397 ( .A(n558), .ZN(n5110) );
  NAND2_X2 U3401 ( .A1(n3151), .A2(n3461), .ZN(n1340) );
  INV_X2 U3404 ( .A(n3193), .ZN(n1341) );
  NAND2_X2 U3405 ( .A1(n3194), .A2(n3160), .ZN(n1342) );
  OAI22_X2 U3406 ( .A1(n5472), .A2(n5360), .B1(n3198), .B2(n3598), .ZN(n5362)
         );
  NAND3_X2 U3407 ( .A1(n3501), .A2(n4525), .A3(n4524), .ZN(n1343) );
  NAND2_X2 U3408 ( .A1(n385), .A2(n1344), .ZN(n3195) );
  INV_X4 U3409 ( .A(n5869), .ZN(n5570) );
  NOR2_X4 U3411 ( .A1(n3772), .A2(n1358), .ZN(n4239) );
  NAND2_X2 U3412 ( .A1(n4218), .A2(n1347), .ZN(n4223) );
  NOR2_X2 U3413 ( .A1(n1349), .A2(n1348), .ZN(n1347) );
  NOR2_X2 U3414 ( .A1(n4216), .A2(n3342), .ZN(n1348) );
  NAND3_X2 U3417 ( .A1(n2127), .A2(n473), .A3(n2899), .ZN(n3585) );
  INV_X4 U3418 ( .A(n4527), .ZN(n2117) );
  NAND2_X4 U3419 ( .A1(n1788), .A2(n1787), .ZN(n1789) );
  NOR2_X2 U3420 ( .A1(n924), .A2(n3143), .ZN(n3159) );
  NOR2_X4 U3423 ( .A1(n2931), .A2(n2775), .ZN(n4577) );
  NAND2_X2 U3424 ( .A1(n1693), .A2(n5794), .ZN(n3353) );
  NAND2_X2 U3426 ( .A1(n3405), .A2(n2603), .ZN(n2605) );
  BUF_X4 U3427 ( .A(n4735), .Z(n1350) );
  NAND2_X2 U3431 ( .A1(n1353), .A2(n1352), .ZN(n1699) );
  NAND2_X2 U3432 ( .A1(n5257), .A2(n3240), .ZN(n1352) );
  NAND2_X2 U3433 ( .A1(n2890), .A2(n5258), .ZN(n1353) );
  INV_X4 U3434 ( .A(n3304), .ZN(n1849) );
  BUF_X4 U3435 ( .A(n606), .Z(n1354) );
  INV_X4 U3436 ( .A(n3326), .ZN(n3242) );
  BUF_X4 U3437 ( .A(n5968), .Z(n1355) );
  INV_X4 U3439 ( .A(n5927), .ZN(n5976) );
  INV_X8 U3440 ( .A(a[21]), .ZN(n1760) );
  NAND2_X4 U3442 ( .A1(n2421), .A2(n2419), .ZN(n1461) );
  NAND2_X2 U3444 ( .A1(n3521), .A2(n3522), .ZN(n1460) );
  NAND3_X2 U3445 ( .A1(n5608), .A2(n2986), .A3(n5607), .ZN(\d[35] ) );
  BUF_X4 U3450 ( .A(n6336), .Z(n1359) );
  NAND2_X2 U3451 ( .A1(n4193), .A2(n4162), .ZN(n2339) );
  NAND2_X2 U3452 ( .A1(n4160), .A2(n4161), .ZN(n4193) );
  NAND2_X2 U3453 ( .A1(n1362), .A2(n986), .ZN(n2566) );
  NAND2_X2 U3454 ( .A1(n4083), .A2(n3702), .ZN(n1363) );
  XOR2_X2 U3455 ( .A(b[6]), .B(a[1]), .Z(n1542) );
  NAND2_X2 U3456 ( .A1(n512), .A2(n184), .ZN(n3327) );
  NAND3_X2 U3457 ( .A1(n1364), .A2(n1365), .A3(n4509), .ZN(n2790) );
  NAND2_X2 U3458 ( .A1(n4508), .A2(n6617), .ZN(n1365) );
  OAI21_X2 U3460 ( .B1(n2803), .B2(n1006), .A(n2144), .ZN(n1572) );
  OAI22_X2 U3461 ( .A1(n568), .A2(b[21]), .B1(n6211), .B2(n5951), .ZN(n2372)
         );
  INV_X2 U3462 ( .A(n2133), .ZN(n2132) );
  NAND3_X2 U3463 ( .A1(n4273), .A2(n2140), .A3(n3462), .ZN(n2133) );
  NAND3_X2 U3464 ( .A1(n5921), .A2(n5919), .A3(n5920), .ZN(n5925) );
  NAND2_X2 U3468 ( .A1(n5780), .A2(n5781), .ZN(n1840) );
  INV_X4 U3469 ( .A(n1841), .ZN(n2375) );
  AOI22_X2 U3470 ( .A1(n1872), .A2(n4452), .B1(n1370), .B2(n1047), .ZN(n4458)
         );
  NOR2_X2 U3472 ( .A1(n440), .A2(n3835), .ZN(n3872) );
  NAND2_X2 U3474 ( .A1(n4941), .A2(n4408), .ZN(n1371) );
  BUF_X4 U3477 ( .A(n4776), .Z(n1765) );
  NOR2_X4 U3478 ( .A1(n1374), .A2(n5383), .ZN(n5622) );
  XNOR2_X1 U3479 ( .A(n6331), .B(n5383), .ZN(n5389) );
  OAI21_X1 U3485 ( .B1(n4914), .B2(n4913), .A(n4915), .ZN(n1381) );
  INV_X8 U3486 ( .A(n5218), .ZN(n5077) );
  NAND3_X4 U3487 ( .A1(n1384), .A2(a[13]), .A3(a[14]), .ZN(n5218) );
  NAND2_X2 U3492 ( .A1(n1387), .A2(n3727), .ZN(n1386) );
  INV_X8 U3493 ( .A(n2098), .ZN(n5190) );
  NAND2_X4 U3494 ( .A1(n1389), .A2(n1388), .ZN(n2098) );
  NAND2_X4 U3495 ( .A1(n2887), .A2(a[21]), .ZN(n1388) );
  INV_X8 U3496 ( .A(a[22]), .ZN(n2887) );
  INV_X8 U3498 ( .A(a[21]), .ZN(n1448) );
  NOR2_X2 U3499 ( .A1(n5187), .A2(n5186), .ZN(n1390) );
  NAND2_X2 U3501 ( .A1(n1393), .A2(n1392), .ZN(n5149) );
  NAND2_X2 U3503 ( .A1(n5077), .A2(b[18]), .ZN(n1393) );
  NOR2_X2 U3504 ( .A1(n5079), .A2(n5078), .ZN(n2489) );
  NAND2_X2 U3505 ( .A1(n5186), .A2(n5187), .ZN(n1394) );
  NAND2_X2 U3507 ( .A1(n5146), .A2(n5145), .ZN(n1395) );
  NOR2_X4 U3508 ( .A1(n1399), .A2(n1396), .ZN(n5186) );
  NAND2_X2 U3509 ( .A1(n1398), .A2(n1397), .ZN(n1396) );
  NAND2_X2 U3510 ( .A1(n2406), .A2(b[17]), .ZN(n1398) );
  NOR2_X4 U3511 ( .A1(n3111), .A2(n5148), .ZN(n1399) );
  XNOR2_X2 U3512 ( .A(n1400), .B(n5757), .ZN(n5763) );
  NAND2_X2 U3513 ( .A1(n1401), .A2(n1402), .ZN(n3474) );
  INV_X2 U3514 ( .A(n3982), .ZN(n1402) );
  NAND2_X2 U3515 ( .A1(n1404), .A2(n1403), .ZN(n3889) );
  INV_X2 U3516 ( .A(n3928), .ZN(n3621) );
  NAND3_X2 U3517 ( .A1(n766), .A2(n1403), .A3(n1050), .ZN(n3928) );
  NOR2_X4 U3519 ( .A1(n395), .A2(a[23]), .ZN(n4752) );
  NAND2_X4 U3520 ( .A1(a[22]), .A2(a[21]), .ZN(n1405) );
  AOI21_X2 U3521 ( .B1(n1407), .B2(n1409), .A(n1411), .ZN(n5263) );
  NAND2_X2 U3523 ( .A1(n5239), .A2(n1036), .ZN(n1409) );
  XNOR2_X2 U3531 ( .A(n1418), .B(n5203), .ZN(n1759) );
  XNOR2_X2 U3532 ( .A(n5152), .B(n5188), .ZN(n5203) );
  NAND2_X2 U3535 ( .A1(n2857), .A2(n2856), .ZN(n5202) );
  NAND2_X2 U3536 ( .A1(n2857), .A2(n2856), .ZN(n1420) );
  AOI21_X2 U3541 ( .B1(n5143), .B2(n5144), .A(n5142), .ZN(n5204) );
  INV_X2 U3542 ( .A(n5153), .ZN(n1425) );
  NOR2_X2 U3543 ( .A1(n1879), .A2(n1878), .ZN(n5153) );
  INV_X4 U3544 ( .A(n1426), .ZN(n5154) );
  NAND2_X2 U3545 ( .A1(n1878), .A2(n1879), .ZN(n1426) );
  NAND2_X2 U3546 ( .A1(n1427), .A2(b[20]), .ZN(n2860) );
  NAND2_X1 U3547 ( .A1(n1427), .A2(b[16]), .ZN(n3374) );
  NAND2_X1 U3548 ( .A1(b[23]), .A2(n1427), .ZN(n2570) );
  NAND2_X2 U3549 ( .A1(n2958), .A2(n6459), .ZN(n1427) );
  NAND2_X2 U3550 ( .A1(n2441), .A2(n1428), .ZN(n5173) );
  NAND3_X2 U3551 ( .A1(n1535), .A2(n1911), .A3(n1910), .ZN(n1430) );
  NAND3_X2 U3552 ( .A1(n1010), .A2(n1514), .A3(n3890), .ZN(n1433) );
  NAND3_X2 U3553 ( .A1(n1433), .A2(n1434), .A3(n1432), .ZN(n1513) );
  INV_X2 U3554 ( .A(n1514), .ZN(n1435) );
  NOR3_X4 U3555 ( .A1(n4607), .A2(n4608), .A3(n4606), .ZN(n4657) );
  INV_X2 U3557 ( .A(n1437), .ZN(n1438) );
  NAND2_X2 U3559 ( .A1(n2549), .A2(n4805), .ZN(n1445) );
  INV_X2 U3560 ( .A(n4808), .ZN(n1446) );
  OAI21_X2 U3561 ( .B1(n1439), .B2(n2030), .A(n341), .ZN(n1443) );
  XNOR2_X2 U3562 ( .A(n4782), .B(n2885), .ZN(n4882) );
  NOR2_X2 U3564 ( .A1(n955), .A2(n1442), .ZN(n1441) );
  NAND3_X2 U3565 ( .A1(n1447), .A2(n1446), .A3(n1445), .ZN(n1444) );
  NOR2_X2 U3566 ( .A1(n1448), .A2(a[20]), .ZN(n3352) );
  BUF_X4 U3567 ( .A(n2283), .Z(n1449) );
  AOI22_X2 U3568 ( .A1(n1998), .A2(n3335), .B1(n1997), .B2(n4585), .ZN(n2283)
         );
  NAND2_X2 U3569 ( .A1(n3554), .A2(n1450), .ZN(n1453) );
  XNOR2_X2 U3570 ( .A(n2545), .B(n4004), .ZN(n3554) );
  OAI21_X2 U3571 ( .B1(n1033), .B2(n2171), .A(n3023), .ZN(n1451) );
  INV_X2 U3572 ( .A(n3023), .ZN(n1454) );
  AOI22_X2 U3573 ( .A1(n2644), .A2(n1456), .B1(n6459), .B2(n4530), .ZN(n1717)
         );
  INV_X2 U3575 ( .A(n4851), .ZN(n4846) );
  NAND2_X2 U3576 ( .A1(n4851), .A2(b[3]), .ZN(n3760) );
  NAND2_X2 U3577 ( .A1(b[3]), .A2(a[23]), .ZN(n4851) );
  INV_X4 U3578 ( .A(n2014), .ZN(n3546) );
  NAND2_X1 U3579 ( .A1(n1640), .A2(n6521), .ZN(n1458) );
  NAND2_X2 U3580 ( .A1(n1460), .A2(n1459), .ZN(n2426) );
  INV_X2 U3581 ( .A(n3523), .ZN(n1459) );
  NAND2_X2 U3582 ( .A1(n1640), .A2(n6521), .ZN(n3522) );
  NAND2_X2 U3584 ( .A1(n6210), .A2(n1461), .ZN(n3567) );
  NAND3_X2 U3586 ( .A1(n1011), .A2(n1055), .A3(n4796), .ZN(n1462) );
  NAND2_X2 U3587 ( .A1(n4799), .A2(n4800), .ZN(n4936) );
  NAND2_X2 U3592 ( .A1(n4717), .A2(n1466), .ZN(n2956) );
  NAND2_X2 U3594 ( .A1(n1469), .A2(n1894), .ZN(n2021) );
  NOR2_X2 U3595 ( .A1(n1985), .A2(n1984), .ZN(n1940) );
  INV_X2 U3596 ( .A(n2613), .ZN(n3467) );
  INV_X2 U3598 ( .A(n1508), .ZN(n1472) );
  INV_X2 U3599 ( .A(n4168), .ZN(n4163) );
  XNOR2_X2 U3600 ( .A(n4164), .B(n4168), .ZN(n2567) );
  AOI22_X2 U3601 ( .A1(n961), .A2(a[0]), .B1(n4219), .B2(n1324), .ZN(n4168) );
  NAND2_X2 U3603 ( .A1(n1474), .A2(n1059), .ZN(n1473) );
  NAND2_X2 U3606 ( .A1(n1479), .A2(n2659), .ZN(n1478) );
  NAND2_X2 U3607 ( .A1(n1481), .A2(n2659), .ZN(n1480) );
  INV_X2 U3608 ( .A(n4937), .ZN(n1481) );
  INV_X2 U3610 ( .A(n4732), .ZN(n1482) );
  AOI21_X1 U3612 ( .B1(n3501), .B2(n4525), .A(n1484), .ZN(n4579) );
  NAND2_X4 U3615 ( .A1(n1657), .A2(n1656), .ZN(n1485) );
  NOR2_X2 U3616 ( .A1(n1486), .A2(n3891), .ZN(n2333) );
  NOR2_X2 U3617 ( .A1(n1487), .A2(n3851), .ZN(n3891) );
  NOR2_X2 U3619 ( .A1(n3617), .A2(n3849), .ZN(n1489) );
  XNOR2_X2 U3620 ( .A(n1491), .B(n3751), .ZN(n2029) );
  NAND2_X2 U3621 ( .A1(n1055), .A2(n4796), .ZN(n1490) );
  NAND2_X2 U3622 ( .A1(n3748), .A2(n1492), .ZN(n1491) );
  OAI21_X2 U3623 ( .B1(n4930), .B2(n4929), .A(n1751), .ZN(n1492) );
  NAND2_X2 U3628 ( .A1(n1495), .A2(n3898), .ZN(n1494) );
  NOR2_X2 U3629 ( .A1(n3897), .A2(n1496), .ZN(n1495) );
  INV_X2 U3630 ( .A(n2277), .ZN(n1496) );
  OAI21_X2 U3631 ( .B1(n1498), .B2(n3897), .A(n3899), .ZN(n1497) );
  NOR2_X2 U3632 ( .A1(n3856), .A2(n3855), .ZN(n3897) );
  NAND2_X2 U3633 ( .A1(n283), .A2(n5321), .ZN(n5767) );
  INV_X4 U3635 ( .A(n1500), .ZN(n2827) );
  INV_X2 U3638 ( .A(n2517), .ZN(n5132) );
  NOR2_X2 U3639 ( .A1(n1505), .A2(n280), .ZN(n5210) );
  NAND2_X2 U3640 ( .A1(n5129), .A2(n5128), .ZN(n5209) );
  NOR2_X2 U3642 ( .A1(n4733), .A2(n3640), .ZN(n1508) );
  XNOR2_X2 U3645 ( .A(n1513), .B(n3895), .ZN(n3860) );
  NOR2_X2 U3646 ( .A1(n1512), .A2(n1511), .ZN(n3895) );
  NAND3_X2 U3647 ( .A1(n1743), .A2(n1741), .A3(n1742), .ZN(n1514) );
  INV_X2 U3649 ( .A(n5004), .ZN(n1516) );
  NAND3_X2 U3650 ( .A1(n415), .A2(n4881), .A3(n2518), .ZN(n1521) );
  NAND2_X4 U3651 ( .A1(n1519), .A2(n1518), .ZN(n4913) );
  NAND2_X2 U3653 ( .A1(n1522), .A2(n1521), .ZN(n4915) );
  NOR2_X4 U3654 ( .A1(n2830), .A2(n4541), .ZN(n1526) );
  NOR2_X2 U3655 ( .A1(n4539), .A2(n4538), .ZN(n1529) );
  NOR2_X2 U3657 ( .A1(n4540), .A2(n3573), .ZN(n1528) );
  OAI22_X2 U3658 ( .A1(n4537), .A2(n6605), .B1(n4536), .B2(n4535), .ZN(n4538)
         );
  BUF_X4 U3659 ( .A(n4910), .Z(n1530) );
  OAI21_X2 U3660 ( .B1(n4893), .B2(n1531), .A(n4892), .ZN(n3197) );
  OAI21_X2 U3661 ( .B1(n3116), .B2(n1864), .A(n1531), .ZN(n3115) );
  NAND2_X2 U3662 ( .A1(n1532), .A2(n5727), .ZN(n3170) );
  NAND2_X2 U3663 ( .A1(n1533), .A2(n2579), .ZN(n1532) );
  NAND2_X2 U3664 ( .A1(n2588), .A2(n5322), .ZN(n1533) );
  INV_X2 U3665 ( .A(n2189), .ZN(n1535) );
  OAI21_X2 U3666 ( .B1(n2707), .B2(n4316), .A(n2951), .ZN(n2588) );
  NAND2_X2 U3670 ( .A1(n4711), .A2(n3222), .ZN(n2682) );
  NAND2_X2 U3671 ( .A1(n3655), .A2(n3862), .ZN(n3938) );
  NAND2_X2 U3672 ( .A1(n3861), .A2(n2100), .ZN(n3862) );
  OAI21_X2 U3673 ( .B1(n2100), .B2(n3861), .A(n3860), .ZN(n3655) );
  AOI21_X2 U3674 ( .B1(n2436), .B2(n3023), .A(n1033), .ZN(n2100) );
  INV_X8 U3675 ( .A(n2524), .ZN(n3598) );
  NAND2_X2 U3676 ( .A1(n3284), .A2(n1546), .ZN(n3645) );
  NAND2_X2 U3679 ( .A1(n4313), .A2(n1548), .ZN(n3534) );
  NAND2_X2 U3680 ( .A1(n2432), .A2(n2431), .ZN(n1550) );
  INV_X2 U3681 ( .A(n2431), .ZN(n1552) );
  NOR2_X4 U3682 ( .A1(n505), .A2(n4821), .ZN(n3431) );
  NAND2_X4 U3683 ( .A1(n3405), .A2(n3993), .ZN(n2432) );
  NOR2_X2 U3684 ( .A1(n1555), .A2(n1817), .ZN(n1561) );
  XNOR2_X2 U3685 ( .A(n1558), .B(n1556), .ZN(n1711) );
  AOI22_X2 U3687 ( .A1(n1870), .A2(n3559), .B1(n1561), .B2(n6209), .ZN(n1560)
         );
  NOR3_X2 U3691 ( .A1(n4344), .A2(n3049), .A3(n3050), .ZN(n2648) );
  OAI21_X2 U3695 ( .B1(n4629), .B2(n4630), .A(n4628), .ZN(n3620) );
  NOR2_X2 U3696 ( .A1(n1572), .A2(n1573), .ZN(n4630) );
  NAND2_X2 U3697 ( .A1(n1712), .A2(n4579), .ZN(n1574) );
  INV_X4 U3698 ( .A(n4580), .ZN(n2608) );
  NAND3_X2 U3699 ( .A1(n6610), .A2(n4404), .A3(n1575), .ZN(n3306) );
  NAND2_X2 U3701 ( .A1(n4403), .A2(n1575), .ZN(n3694) );
  INV_X2 U3702 ( .A(n1575), .ZN(n4402) );
  NOR2_X2 U3704 ( .A1(n1579), .A2(n4760), .ZN(n1577) );
  INV_X2 U3705 ( .A(n1580), .ZN(n1579) );
  OAI22_X2 U3706 ( .A1(n4690), .A2(n6605), .B1(n4948), .B2(n3683), .ZN(n4692)
         );
  NOR2_X2 U3707 ( .A1(n4693), .A2(n2700), .ZN(n3404) );
  NAND2_X2 U3708 ( .A1(n1028), .A2(n2804), .ZN(n4643) );
  NAND4_X1 U3709 ( .A1(n324), .A2(n1581), .A3(n1028), .A4(n2804), .ZN(n2150)
         );
  NAND3_X2 U3710 ( .A1(n2712), .A2(n511), .A3(n2806), .ZN(n2804) );
  NAND2_X2 U3711 ( .A1(n1949), .A2(n46), .ZN(n1584) );
  NAND2_X2 U3713 ( .A1(n1588), .A2(n1589), .ZN(n1587) );
  INV_X2 U3714 ( .A(n1590), .ZN(n1589) );
  INV_X4 U3715 ( .A(n2322), .ZN(n2443) );
  AOI21_X2 U3718 ( .B1(n3898), .B2(n3899), .A(n3897), .ZN(n3936) );
  NAND2_X2 U3720 ( .A1(n1594), .A2(n3125), .ZN(n1596) );
  NAND2_X2 U3721 ( .A1(n1596), .A2(n1595), .ZN(n5789) );
  OAI21_X2 U3723 ( .B1(n1598), .B2(n2601), .A(n1597), .ZN(n2087) );
  NAND2_X1 U3724 ( .A1(n1599), .A2(n4582), .ZN(n1597) );
  NAND3_X4 U3726 ( .A1(n1760), .A2(a[19]), .A3(a[20]), .ZN(n5895) );
  NOR2_X2 U3727 ( .A1(n369), .A2(n5999), .ZN(n5932) );
  OAI21_X2 U3728 ( .B1(n1604), .B2(n6078), .A(n2332), .ZN(n2331) );
  AOI22_X2 U3729 ( .A1(n1607), .A2(n1605), .B1(n5931), .B2(n1020), .ZN(n1604)
         );
  NOR2_X2 U3730 ( .A1(n369), .A2(n1606), .ZN(n1605) );
  INV_X2 U3731 ( .A(n1020), .ZN(n1606) );
  NAND2_X2 U3732 ( .A1(n1614), .A2(n1613), .ZN(n5489) );
  XNOR2_X2 U3733 ( .A(n5488), .B(n5487), .ZN(n1612) );
  NAND3_X2 U3734 ( .A1(n5434), .A2(n5433), .A3(n1616), .ZN(n1613) );
  INV_X2 U3735 ( .A(n1615), .ZN(n1614) );
  AOI21_X2 U3736 ( .B1(n5434), .B2(n5433), .A(n1616), .ZN(n1615) );
  INV_X2 U3737 ( .A(n5435), .ZN(n1616) );
  AOI21_X2 U3738 ( .B1(n5465), .B2(n5464), .A(n5463), .ZN(n5488) );
  INV_X2 U3739 ( .A(n3548), .ZN(n3549) );
  NAND3_X2 U3740 ( .A1(n1618), .A2(n1617), .A3(n970), .ZN(n3548) );
  NAND2_X2 U3741 ( .A1(n2514), .A2(b[20]), .ZN(n1617) );
  NAND2_X2 U3745 ( .A1(n5009), .A2(n5010), .ZN(n1624) );
  AOI22_X2 U3746 ( .A1(n4088), .A2(n4102), .B1(n1052), .B2(n4100), .ZN(n1626)
         );
  OAI21_X2 U3747 ( .B1(n5214), .B2(n1627), .A(n5213), .ZN(n5598) );
  NAND2_X2 U3748 ( .A1(n1629), .A2(n5177), .ZN(n1631) );
  NOR2_X2 U3752 ( .A1(n1637), .A2(n5091), .ZN(n1745) );
  INV_X2 U3753 ( .A(n3379), .ZN(n1635) );
  NAND3_X2 U3754 ( .A1(n6451), .A2(n5088), .A3(n2799), .ZN(n1638) );
  NOR2_X2 U3755 ( .A1(n2798), .A2(n2797), .ZN(n1639) );
  NAND2_X2 U3756 ( .A1(n1642), .A2(n3382), .ZN(n2417) );
  OAI21_X2 U3759 ( .B1(n1643), .B2(n4859), .A(n2888), .ZN(n2191) );
  NAND2_X2 U3760 ( .A1(n2193), .A2(n2192), .ZN(n1643) );
  NAND2_X2 U3763 ( .A1(n1645), .A2(n3243), .ZN(n4515) );
  NAND2_X2 U3764 ( .A1(b[23]), .A2(n3137), .ZN(n1647) );
  NOR2_X4 U3766 ( .A1(n1652), .A2(n4594), .ZN(n3752) );
  NOR2_X4 U3767 ( .A1(n4592), .A2(n4591), .ZN(n1652) );
  NAND2_X2 U3768 ( .A1(n1846), .A2(n1845), .ZN(n2488) );
  INV_X2 U3769 ( .A(n5038), .ZN(n1655) );
  NAND2_X2 U3771 ( .A1(n1658), .A2(n3107), .ZN(n1656) );
  NAND2_X2 U3772 ( .A1(n567), .A2(n60), .ZN(n1657) );
  BUF_X4 U3773 ( .A(n4892), .Z(n1659) );
  NAND2_X2 U3774 ( .A1(n4880), .A2(n2827), .ZN(n4893) );
  XNOR2_X2 U3776 ( .A(n2837), .B(n1022), .ZN(n1667) );
  XNOR2_X2 U3777 ( .A(n1668), .B(n5890), .ZN(n5545) );
  NOR2_X2 U3778 ( .A1(n1669), .A2(n5891), .ZN(n1668) );
  NOR2_X2 U3779 ( .A1(n5534), .A2(n5533), .ZN(n5891) );
  INV_X2 U3780 ( .A(n5889), .ZN(n1669) );
  NAND2_X2 U3781 ( .A1(n5534), .A2(n5533), .ZN(n5889) );
  AOI21_X2 U3784 ( .B1(n1671), .B2(n1670), .A(n4773), .ZN(n4803) );
  NAND2_X2 U3785 ( .A1(n3242), .A2(n3438), .ZN(n1670) );
  NAND2_X2 U3786 ( .A1(n4772), .A2(b[19]), .ZN(n1671) );
  NOR2_X4 U3788 ( .A1(a[19]), .A2(a[21]), .ZN(n1674) );
  NAND3_X2 U3789 ( .A1(n5916), .A2(n1675), .A3(n5915), .ZN(n5917) );
  NOR3_X2 U3790 ( .A1(n6074), .A2(n5914), .A3(n5913), .ZN(n1675) );
  NAND2_X2 U3791 ( .A1(n1677), .A2(n1676), .ZN(n5893) );
  NAND2_X2 U3792 ( .A1(n1680), .A2(n1679), .ZN(n1677) );
  NOR2_X2 U3794 ( .A1(n3270), .A2(n5411), .ZN(n1680) );
  BUF_X4 U3795 ( .A(n2469), .Z(n1682) );
  NAND2_X2 U3798 ( .A1(n1687), .A2(n1686), .ZN(n4268) );
  NAND2_X2 U3799 ( .A1(n2326), .A2(n3830), .ZN(n4269) );
  INV_X2 U3800 ( .A(n4268), .ZN(n1688) );
  OAI21_X2 U3801 ( .B1(n3353), .B2(n3428), .A(n274), .ZN(n3321) );
  NAND2_X2 U3802 ( .A1(n6206), .A2(n4972), .ZN(n2903) );
  AOI21_X2 U3803 ( .B1(n290), .B2(n3168), .A(n2681), .ZN(n4972) );
  NAND2_X2 U3804 ( .A1(n2268), .A2(n2267), .ZN(n2266) );
  NOR2_X2 U3807 ( .A1(n1695), .A2(n1694), .ZN(n1693) );
  NAND2_X2 U3808 ( .A1(n2637), .A2(n3625), .ZN(n1695) );
  NAND3_X2 U3809 ( .A1(n5629), .A2(n5630), .A3(n1697), .ZN(n2955) );
  NAND2_X2 U3810 ( .A1(n2398), .A2(n5317), .ZN(n1697) );
  AOI22_X2 U3811 ( .A1(n2891), .A2(n1023), .B1(n5331), .B2(n5332), .ZN(n1698)
         );
  NAND2_X2 U3812 ( .A1(n1699), .A2(n5207), .ZN(n5216) );
  NOR2_X2 U3813 ( .A1(n1699), .A2(n5207), .ZN(n5206) );
  NAND3_X2 U3814 ( .A1(n5261), .A2(n5307), .A3(n5262), .ZN(n1701) );
  NAND2_X2 U3815 ( .A1(n5309), .A2(n1001), .ZN(n1702) );
  NAND3_X2 U3817 ( .A1(n4700), .A2(n733), .A3(n4821), .ZN(n1703) );
  INV_X2 U3818 ( .A(n4702), .ZN(n1704) );
  AOI22_X2 U3819 ( .A1(n4698), .A2(a[4]), .B1(n1706), .B2(n1066), .ZN(n1705)
         );
  NAND2_X2 U3820 ( .A1(n1708), .A2(n1707), .ZN(n1706) );
  NAND2_X2 U3821 ( .A1(b[21]), .A2(n733), .ZN(n1707) );
  NAND2_X2 U3822 ( .A1(n566), .A2(n4821), .ZN(n1708) );
  OAI22_X2 U3824 ( .A1(n2830), .A2(n4419), .B1(n4420), .B2(n4421), .ZN(n1710)
         );
  NAND2_X1 U3825 ( .A1(n1711), .A2(n3314), .ZN(n2624) );
  NAND2_X4 U3826 ( .A1(n1713), .A2(n4978), .ZN(n4976) );
  NAND2_X2 U3827 ( .A1(n1530), .A2(n6520), .ZN(n4978) );
  INV_X1 U3828 ( .A(n4899), .ZN(n1715) );
  INV_X2 U3830 ( .A(n2942), .ZN(n1718) );
  NAND2_X2 U3831 ( .A1(n4584), .A2(n2947), .ZN(n2942) );
  NAND2_X4 U3832 ( .A1(n2998), .A2(n3712), .ZN(n4584) );
  NAND2_X2 U3833 ( .A1(n1722), .A2(n1719), .ZN(n2861) );
  INV_X2 U3834 ( .A(n5353), .ZN(n1720) );
  INV_X2 U3835 ( .A(n1723), .ZN(n1722) );
  XNOR2_X2 U3836 ( .A(n2062), .B(n5490), .ZN(n5564) );
  NAND2_X2 U3837 ( .A1(n2063), .A2(n5353), .ZN(n5566) );
  XNOR2_X2 U3838 ( .A(n1724), .B(n5556), .ZN(n5565) );
  NOR2_X2 U3839 ( .A1(n2595), .A2(n4789), .ZN(n1725) );
  AOI21_X2 U3840 ( .B1(n2656), .B2(n5293), .A(n4787), .ZN(n2595) );
  INV_X2 U3841 ( .A(n2596), .ZN(n1726) );
  NAND2_X2 U3844 ( .A1(n1732), .A2(n1731), .ZN(n1730) );
  INV_X2 U3845 ( .A(n5296), .ZN(n1731) );
  INV_X4 U3846 ( .A(n2757), .ZN(n3107) );
  NOR2_X2 U3847 ( .A1(n4405), .A2(n3572), .ZN(n1734) );
  NAND2_X2 U3848 ( .A1(n1738), .A2(n1737), .ZN(n1736) );
  NAND2_X2 U3849 ( .A1(n2656), .A2(b[1]), .ZN(n1740) );
  NAND3_X1 U3851 ( .A1(n2958), .A2(b[1]), .A3(n6459), .ZN(n1743) );
  INV_X2 U3852 ( .A(n1888), .ZN(n3402) );
  NAND2_X2 U3854 ( .A1(n4922), .A2(n6459), .ZN(n1888) );
  NOR2_X2 U3855 ( .A1(n5154), .A2(n5153), .ZN(n1746) );
  AOI21_X2 U3856 ( .B1(n759), .B2(n3108), .A(n6330), .ZN(n1748) );
  AOI21_X2 U3858 ( .B1(n4477), .B2(n4478), .A(n1841), .ZN(n1754) );
  NAND2_X2 U3859 ( .A1(n2367), .A2(n2365), .ZN(n4479) );
  NAND2_X2 U3860 ( .A1(n1754), .A2(n4479), .ZN(n1752) );
  NAND3_X2 U3861 ( .A1(n539), .A2(n6149), .A3(n4472), .ZN(n1755) );
  INV_X4 U3862 ( .A(n1757), .ZN(n4937) );
  NAND2_X4 U3863 ( .A1(n1758), .A2(n4937), .ZN(n3106) );
  NAND2_X1 U3866 ( .A1(n1759), .A2(n821), .ZN(n5213) );
  NOR2_X1 U3867 ( .A1(n1759), .A2(n821), .ZN(n5214) );
  NOR3_X4 U3868 ( .A1(n4989), .A2(a[19]), .A3(a[20]), .ZN(n1763) );
  BUF_X4 U3869 ( .A(n5473), .Z(n1761) );
  BUF_X4 U3870 ( .A(n5473), .Z(n1762) );
  INV_X8 U3871 ( .A(n1763), .ZN(n5473) );
  NOR2_X2 U3875 ( .A1(n1768), .A2(n1767), .ZN(n1766) );
  NAND2_X2 U3876 ( .A1(n6619), .A2(n2279), .ZN(n1769) );
  INV_X2 U3877 ( .A(n1769), .ZN(n1996) );
  XNOR2_X2 U3880 ( .A(n4116), .B(n4114), .ZN(n1771) );
  NAND2_X2 U3882 ( .A1(n4109), .A2(n1773), .ZN(n4116) );
  NOR2_X2 U3883 ( .A1(n4216), .A2(n3538), .ZN(n1774) );
  INV_X2 U3888 ( .A(n2273), .ZN(n1778) );
  NAND2_X2 U3890 ( .A1(n3538), .A2(n1308), .ZN(n4208) );
  NAND2_X2 U3891 ( .A1(n4082), .A2(n1847), .ZN(n2335) );
  NAND2_X4 U3892 ( .A1(n3877), .A2(a[7]), .ZN(n1847) );
  NAND2_X2 U3893 ( .A1(n1779), .A2(n1782), .ZN(n1805) );
  NAND2_X2 U3894 ( .A1(n2352), .A2(n3449), .ZN(n1783) );
  OAI22_X2 U3897 ( .A1(n4757), .A2(n4756), .B1(n4755), .B2(n1455), .ZN(n4865)
         );
  NAND2_X2 U3898 ( .A1(n4759), .A2(n4758), .ZN(n1787) );
  AOI22_X2 U3899 ( .A1(b[9]), .A2(n2382), .B1(n2510), .B2(n6221), .ZN(n4710)
         );
  NOR2_X2 U3901 ( .A1(n1793), .A2(n1792), .ZN(n4758) );
  NAND2_X2 U3904 ( .A1(n1795), .A2(n4859), .ZN(n2190) );
  NOR2_X2 U3905 ( .A1(n1801), .A2(n1803), .ZN(n2590) );
  NAND3_X2 U3907 ( .A1(n1797), .A2(n5019), .A3(n1796), .ZN(n5062) );
  NAND3_X2 U3908 ( .A1(n1802), .A2(n5018), .A3(n1803), .ZN(n1796) );
  NAND3_X2 U3909 ( .A1(n5018), .A2(n1802), .A3(n1801), .ZN(n1797) );
  INV_X2 U3911 ( .A(n5016), .ZN(n1802) );
  INV_X2 U3912 ( .A(n1875), .ZN(n1816) );
  INV_X2 U3913 ( .A(n1815), .ZN(n1813) );
  NAND2_X2 U3916 ( .A1(n1809), .A2(n1806), .ZN(n1878) );
  NAND2_X2 U3919 ( .A1(n6303), .A2(n1814), .ZN(n1809) );
  NAND2_X2 U3921 ( .A1(n1812), .A2(n1811), .ZN(n1879) );
  NAND3_X2 U3922 ( .A1(n1032), .A2(n1816), .A3(n1815), .ZN(n1811) );
  BUF_X4 U3924 ( .A(n3232), .Z(n1818) );
  NOR2_X4 U3925 ( .A1(n1821), .A2(n1819), .ZN(n2033) );
  NOR2_X2 U3926 ( .A1(n1822), .A2(n1818), .ZN(n1819) );
  AOI21_X2 U3927 ( .B1(n1822), .B2(n1818), .A(n538), .ZN(n1821) );
  AOI22_X2 U3929 ( .A1(b[1]), .A2(n3581), .B1(n1326), .B2(n1823), .ZN(n1825)
         );
  NOR2_X2 U3936 ( .A1(n1831), .A2(n629), .ZN(n3076) );
  NAND2_X2 U3937 ( .A1(n2990), .A2(n3229), .ZN(n1834) );
  OAI22_X2 U3941 ( .A1(n5079), .A2(n4052), .B1(n4053), .B2(n4054), .ZN(n1838)
         );
  OAI21_X2 U3943 ( .B1(n4465), .B2(n4464), .A(n4463), .ZN(n4478) );
  NAND2_X2 U3944 ( .A1(n1842), .A2(n1843), .ZN(n4477) );
  NAND2_X2 U3945 ( .A1(n4069), .A2(n4068), .ZN(n4463) );
  NAND2_X1 U3948 ( .A1(n2765), .A2(n6329), .ZN(n1951) );
  OAI21_X2 U3950 ( .B1(n1857), .B2(n1856), .A(n1855), .ZN(n1854) );
  NOR2_X2 U3952 ( .A1(n3752), .A2(n2825), .ZN(n1856) );
  NAND2_X2 U3953 ( .A1(n1859), .A2(n1858), .ZN(n4671) );
  NAND2_X2 U3954 ( .A1(n1861), .A2(n1860), .ZN(n1859) );
  INV_X1 U3955 ( .A(n3268), .ZN(n1860) );
  NAND2_X2 U3956 ( .A1(n3291), .A2(n3290), .ZN(n1861) );
  INV_X2 U3957 ( .A(n1659), .ZN(n1862) );
  NAND2_X2 U3958 ( .A1(n987), .A2(n3115), .ZN(n1863) );
  XNOR2_X2 U3959 ( .A(n1865), .B(n4001), .ZN(n2544) );
  NAND2_X2 U3961 ( .A1(n3169), .A2(n3168), .ZN(n2895) );
  AOI22_X2 U3962 ( .A1(n2033), .A2(n1866), .B1(n641), .B2(n2708), .ZN(n3168)
         );
  NAND2_X2 U3964 ( .A1(n1868), .A2(n5789), .ZN(n3169) );
  NAND2_X2 U3965 ( .A1(n6602), .A2(n2034), .ZN(n1868) );
  INV_X1 U3967 ( .A(n1870), .ZN(n3314) );
  NAND2_X2 U3968 ( .A1(n5001), .A2(n5000), .ZN(n5052) );
  NAND2_X2 U3969 ( .A1(n4451), .A2(n1873), .ZN(n1872) );
  NOR2_X2 U3970 ( .A1(n5122), .A2(n5123), .ZN(n1875) );
  NAND2_X2 U3971 ( .A1(n2356), .A2(n2355), .ZN(n5123) );
  NAND2_X2 U3974 ( .A1(n3574), .A2(n432), .ZN(n3093) );
  XNOR2_X2 U3975 ( .A(n5296), .B(n5294), .ZN(n1877) );
  NAND3_X2 U3976 ( .A1(n3429), .A2(n4551), .A3(n3510), .ZN(n1881) );
  INV_X2 U3977 ( .A(n4236), .ZN(n3358) );
  NOR2_X2 U3978 ( .A1(n4236), .A2(n1884), .ZN(n1883) );
  NAND2_X2 U3982 ( .A1(n3312), .A2(n6263), .ZN(n1936) );
  INV_X4 U3984 ( .A(n1889), .ZN(n5174) );
  NAND2_X2 U3985 ( .A1(n1890), .A2(n5175), .ZN(n2857) );
  NAND2_X2 U3986 ( .A1(n5174), .A2(n5173), .ZN(n1890) );
  XNOR2_X2 U3987 ( .A(n4036), .B(n4035), .ZN(n1891) );
  AOI21_X2 U3988 ( .B1(n6459), .B2(n3956), .A(n3955), .ZN(n4036) );
  NAND3_X2 U3989 ( .A1(n4043), .A2(n4042), .A3(n4040), .ZN(n1892) );
  NAND2_X2 U3990 ( .A1(n1894), .A2(n2003), .ZN(n2002) );
  NAND2_X2 U3991 ( .A1(n1895), .A2(n3540), .ZN(n4560) );
  INV_X2 U3993 ( .A(n4812), .ZN(n1895) );
  XNOR2_X1 U3994 ( .A(n4812), .B(n1896), .ZN(n6104) );
  NAND2_X2 U3996 ( .A1(n4255), .A2(n4287), .ZN(n1899) );
  NAND2_X2 U3997 ( .A1(n4253), .A2(n4254), .ZN(n4287) );
  INV_X1 U4001 ( .A(n1902), .ZN(n2320) );
  NOR2_X1 U4003 ( .A1(n6009), .A2(n1902), .ZN(n3612) );
  NAND2_X1 U4004 ( .A1(n5974), .A2(n1902), .ZN(n5979) );
  NAND2_X2 U4005 ( .A1(n1903), .A2(n1905), .ZN(n4979) );
  NAND2_X2 U4006 ( .A1(n1904), .A2(n891), .ZN(n1903) );
  NAND2_X2 U4007 ( .A1(n1907), .A2(n1906), .ZN(n1905) );
  AOI22_X2 U4008 ( .A1(n2677), .A2(n5092), .B1(n3093), .B2(n3341), .ZN(n1906)
         );
  NAND2_X2 U4009 ( .A1(n2884), .A2(n2883), .ZN(n3341) );
  NOR2_X2 U4011 ( .A1(n2549), .A2(n4805), .ZN(n2030) );
  INV_X2 U4013 ( .A(n3862), .ZN(n1912) );
  XNOR2_X2 U4014 ( .A(n2649), .B(n3886), .ZN(n3654) );
  XNOR2_X1 U4016 ( .A(n6381), .B(n5662), .ZN(n5663) );
  INV_X8 U4017 ( .A(a[13]), .ZN(n1916) );
  NOR2_X2 U4019 ( .A1(n1922), .A2(n3812), .ZN(n2171) );
  NAND3_X2 U4020 ( .A1(n3997), .A2(n2432), .A3(n2431), .ZN(n4247) );
  BUF_X4 U4022 ( .A(n3711), .Z(n1923) );
  NAND3_X2 U4023 ( .A1(n1923), .A2(n1926), .A3(n2470), .ZN(n1924) );
  NAND2_X2 U4028 ( .A1(n1931), .A2(n1930), .ZN(n4566) );
  INV_X2 U4029 ( .A(n3577), .ZN(n1931) );
  INV_X4 U4030 ( .A(n4940), .ZN(n5109) );
  AOI22_X2 U4033 ( .A1(n1936), .A2(n5022), .B1(n6460), .B2(b[7]), .ZN(n5064)
         );
  NAND2_X2 U4034 ( .A1(n1937), .A2(n4684), .ZN(n4717) );
  NAND2_X2 U4035 ( .A1(n1939), .A2(n1938), .ZN(n1937) );
  NAND2_X4 U4037 ( .A1(a[8]), .A2(a[7]), .ZN(n4998) );
  INV_X2 U4038 ( .A(n4573), .ZN(n4572) );
  NAND2_X2 U4040 ( .A1(n1183), .A2(n3074), .ZN(n5040) );
  NAND2_X2 U4043 ( .A1(n891), .A2(n3370), .ZN(n1946) );
  NAND2_X2 U4045 ( .A1(n4874), .A2(n1949), .ZN(n4875) );
  INV_X2 U4047 ( .A(n2680), .ZN(n1950) );
  NAND2_X2 U4049 ( .A1(n1831), .A2(n4959), .ZN(n1954) );
  INV_X2 U4050 ( .A(n4838), .ZN(n1956) );
  NAND2_X2 U4051 ( .A1(n1959), .A2(n1958), .ZN(n2350) );
  NAND3_X2 U4052 ( .A1(n1960), .A2(n2399), .A3(n4744), .ZN(n1958) );
  NAND3_X2 U4053 ( .A1(n5132), .A2(n1031), .A3(n5130), .ZN(n3109) );
  NAND2_X2 U4056 ( .A1(n1963), .A2(n1961), .ZN(n4079) );
  INV_X2 U4057 ( .A(n4077), .ZN(n1962) );
  INV_X2 U4058 ( .A(n4075), .ZN(n1964) );
  NAND2_X2 U4061 ( .A1(n1967), .A2(n1966), .ZN(n1965) );
  INV_X2 U4062 ( .A(n3747), .ZN(n1966) );
  NAND2_X2 U4063 ( .A1(n1038), .A2(n1970), .ZN(n1967) );
  NAND3_X2 U4064 ( .A1(n1970), .A2(n1038), .A3(n3747), .ZN(n1968) );
  NAND2_X2 U4067 ( .A1(n3965), .A2(n6251), .ZN(n1970) );
  OAI21_X2 U4068 ( .B1(n5079), .B2(n3925), .A(n2996), .ZN(n3965) );
  INV_X2 U4070 ( .A(n5048), .ZN(n2764) );
  NOR2_X2 U4071 ( .A1(n3630), .A2(n3631), .ZN(n5048) );
  NAND2_X2 U4072 ( .A1(n2116), .A2(n2115), .ZN(n3630) );
  NAND2_X1 U4073 ( .A1(n189), .A2(n1973), .ZN(n3216) );
  NAND2_X2 U4075 ( .A1(n1976), .A2(n3078), .ZN(n3079) );
  NOR2_X2 U4076 ( .A1(n2577), .A2(a[14]), .ZN(n4415) );
  INV_X8 U4078 ( .A(n5219), .ZN(n5076) );
  NAND2_X2 U4082 ( .A1(n3385), .A2(n3251), .ZN(n1989) );
  NAND2_X2 U4083 ( .A1(n1994), .A2(n1993), .ZN(n1992) );
  NAND2_X2 U4085 ( .A1(n2947), .A2(n4584), .ZN(n1998) );
  NAND2_X2 U4086 ( .A1(n2727), .A2(n1999), .ZN(n2472) );
  NAND2_X2 U4088 ( .A1(n4745), .A2(n1999), .ZN(n4836) );
  NAND2_X1 U4089 ( .A1(n4949), .A2(n1999), .ZN(n4950) );
  AOI22_X2 U4090 ( .A1(n3908), .A2(n3907), .B1(n3906), .B2(n1999), .ZN(n3942)
         );
  NOR2_X1 U4092 ( .A1(n4417), .A2(n6588), .ZN(n2000) );
  NAND2_X4 U4095 ( .A1(n2002), .A2(n6357), .ZN(n5859) );
  AOI22_X2 U4097 ( .A1(n5326), .A2(n1016), .B1(n2154), .B2(n5325), .ZN(n5327)
         );
  OAI21_X2 U4099 ( .B1(n4644), .B2(n4528), .A(n4639), .ZN(n5834) );
  NAND2_X2 U4100 ( .A1(n2008), .A2(n5794), .ZN(n2007) );
  NAND2_X2 U4101 ( .A1(n3626), .A2(n3940), .ZN(n2531) );
  NAND2_X2 U4105 ( .A1(n3152), .A2(n3304), .ZN(n2014) );
  NAND2_X2 U4106 ( .A1(n4503), .A2(n3439), .ZN(n4551) );
  NAND2_X4 U4107 ( .A1(n3510), .A2(n4550), .ZN(n4552) );
  INV_X2 U4108 ( .A(n4638), .ZN(n2267) );
  OAI21_X2 U4109 ( .B1(n2016), .B2(n2015), .A(n4081), .ZN(n4638) );
  NOR2_X2 U4110 ( .A1(n4080), .A2(n4079), .ZN(n2015) );
  INV_X8 U4112 ( .A(n3729), .ZN(n4405) );
  NAND3_X2 U4113 ( .A1(b[21]), .A2(n4492), .A3(n1064), .ZN(n4493) );
  NOR2_X2 U4114 ( .A1(n4588), .A2(n1064), .ZN(n4659) );
  AOI21_X1 U4115 ( .B1(n4129), .B2(n1064), .A(n4492), .ZN(n4133) );
  NAND2_X2 U4117 ( .A1(n2582), .A2(n2446), .ZN(n2020) );
  NAND2_X2 U4118 ( .A1(n2632), .A2(n2631), .ZN(n2027) );
  INV_X1 U4119 ( .A(n4731), .ZN(n2630) );
  NAND2_X2 U4120 ( .A1(n2251), .A2(n2254), .ZN(n4808) );
  XNOR2_X2 U4121 ( .A(n4568), .B(n4567), .ZN(n2031) );
  INV_X8 U4122 ( .A(a[19]), .ZN(n2032) );
  OAI22_X2 U4123 ( .A1(n3326), .A2(b[17]), .B1(n3217), .B2(n3581), .ZN(n2035)
         );
  NOR2_X2 U4124 ( .A1(n2801), .A2(n2800), .ZN(n4732) );
  NOR2_X4 U4126 ( .A1(a[21]), .A2(a[22]), .ZN(n2038) );
  NAND2_X2 U4127 ( .A1(n4191), .A2(n4190), .ZN(n2376) );
  INV_X2 U4129 ( .A(n2041), .ZN(n3255) );
  NAND2_X2 U4132 ( .A1(n808), .A2(n5012), .ZN(n3669) );
  NAND2_X4 U4133 ( .A1(a[16]), .A2(a[15]), .ZN(n2045) );
  INV_X4 U4134 ( .A(n3532), .ZN(n2047) );
  INV_X2 U4136 ( .A(n3531), .ZN(n2046) );
  NAND2_X2 U4137 ( .A1(n5081), .A2(n5082), .ZN(n2050) );
  NOR2_X4 U4138 ( .A1(n3531), .A2(n3532), .ZN(n5081) );
  XNOR2_X2 U4142 ( .A(n5368), .B(n2814), .ZN(n2813) );
  NAND3_X2 U4143 ( .A1(n2053), .A2(n3599), .A3(n2052), .ZN(n2814) );
  NAND2_X2 U4144 ( .A1(n2514), .A2(b[16]), .ZN(n2052) );
  NAND2_X2 U4145 ( .A1(n2055), .A2(n2817), .ZN(n2054) );
  NAND2_X2 U4146 ( .A1(n2058), .A2(n2057), .ZN(n4805) );
  NAND2_X2 U4147 ( .A1(n2739), .A2(n3562), .ZN(n2057) );
  NOR2_X2 U4149 ( .A1(n2059), .A2(n5371), .ZN(n5875) );
  NAND2_X2 U4150 ( .A1(n5290), .A2(n6150), .ZN(n2060) );
  NAND2_X2 U4151 ( .A1(n3558), .A2(n6152), .ZN(n2061) );
  NOR2_X2 U4152 ( .A1(n5492), .A2(n5491), .ZN(n2062) );
  NAND2_X2 U4155 ( .A1(n2067), .A2(n5567), .ZN(n5610) );
  NAND2_X2 U4157 ( .A1(n2069), .A2(n2068), .ZN(n2071) );
  NAND2_X2 U4159 ( .A1(n2071), .A2(n2070), .ZN(n5514) );
  NAND4_X1 U4160 ( .A1(n972), .A2(n5502), .A3(n5508), .A4(n5503), .ZN(n2070)
         );
  NOR2_X2 U4161 ( .A1(n5514), .A2(n5513), .ZN(n2072) );
  NAND2_X2 U4163 ( .A1(n3028), .A2(n3027), .ZN(n2073) );
  OAI22_X2 U4165 ( .A1(n2076), .A2(n2075), .B1(n5114), .B2(n5113), .ZN(n5116)
         );
  NOR2_X2 U4166 ( .A1(n3449), .A2(n5112), .ZN(n2075) );
  NAND2_X2 U4167 ( .A1(n3308), .A2(n4996), .ZN(n5083) );
  NAND2_X2 U4169 ( .A1(n2078), .A2(n2077), .ZN(n5195) );
  NAND2_X2 U4170 ( .A1(n3230), .A2(n5293), .ZN(n2078) );
  NAND2_X1 U4171 ( .A1(n3189), .A2(n3188), .ZN(n2079) );
  BUF_X4 U4172 ( .A(n2087), .Z(n2086) );
  INV_X2 U4173 ( .A(n3569), .ZN(n2088) );
  NAND2_X1 U4177 ( .A1(n2335), .A2(n2095), .ZN(n4162) );
  INV_X8 U4178 ( .A(n4491), .ZN(n4219) );
  BUF_X4 U4179 ( .A(n2100), .Z(n2099) );
  INV_X4 U4180 ( .A(n4581), .ZN(n2102) );
  NAND2_X2 U4181 ( .A1(n2101), .A2(n4581), .ZN(n2691) );
  NAND2_X2 U4182 ( .A1(n2103), .A2(b[0]), .ZN(n2104) );
  NAND2_X2 U4183 ( .A1(n6344), .A2(n3674), .ZN(n3239) );
  OAI21_X2 U4184 ( .B1(n3347), .B2(n3060), .A(n4470), .ZN(n3674) );
  NAND2_X2 U4185 ( .A1(n2105), .A2(n2106), .ZN(n3266) );
  NAND3_X2 U4186 ( .A1(n2317), .A2(n486), .A3(n2774), .ZN(n2105) );
  INV_X2 U4187 ( .A(n2108), .ZN(n5142) );
  NAND2_X2 U4188 ( .A1(n2761), .A2(n2763), .ZN(n2108) );
  NAND3_X2 U4189 ( .A1(n2112), .A2(n485), .A3(n3174), .ZN(n3981) );
  NAND2_X2 U4190 ( .A1(n4278), .A2(n4277), .ZN(n2113) );
  NOR2_X2 U4192 ( .A1(n2428), .A2(n2429), .ZN(n4281) );
  NAND2_X2 U4193 ( .A1(n2675), .A2(b[21]), .ZN(n2115) );
  INV_X8 U4195 ( .A(n4886), .ZN(n5074) );
  NAND2_X2 U4196 ( .A1(n2123), .A2(n2121), .ZN(n3730) );
  NAND2_X1 U4197 ( .A1(n2326), .A2(n4326), .ZN(n2123) );
  NAND2_X2 U4198 ( .A1(n3739), .A2(n3740), .ZN(n4322) );
  INV_X4 U4199 ( .A(n2681), .ZN(n2127) );
  NOR2_X4 U4200 ( .A1(n3671), .A2(a[3]), .ZN(n3729) );
  NOR2_X4 U4201 ( .A1(a[1]), .A2(a[2]), .ZN(n4677) );
  INV_X2 U4202 ( .A(n2131), .ZN(n4339) );
  INV_X2 U4205 ( .A(n2139), .ZN(n2138) );
  NAND2_X2 U4208 ( .A1(n2143), .A2(n6155), .ZN(n2142) );
  NAND2_X2 U4211 ( .A1(n2804), .A2(n1028), .ZN(n2149) );
  OAI21_X2 U4213 ( .B1(n4973), .B2(n4974), .A(n5919), .ZN(n3407) );
  AOI21_X2 U4215 ( .B1(n2676), .B2(n4325), .A(n2158), .ZN(n3051) );
  NAND2_X2 U4216 ( .A1(n2159), .A2(n2402), .ZN(n2158) );
  NAND2_X2 U4217 ( .A1(n2160), .A2(n4322), .ZN(n2402) );
  AOI21_X2 U4218 ( .B1(n1762), .B2(b[1]), .A(n4324), .ZN(n4435) );
  INV_X8 U4220 ( .A(a[7]), .ZN(n2162) );
  INV_X2 U4221 ( .A(n4632), .ZN(n2667) );
  OAI22_X2 U4222 ( .A1(n2165), .A2(n4642), .B1(n4646), .B2(n2164), .ZN(n4632)
         );
  NOR2_X2 U4223 ( .A1(n4557), .A2(n4643), .ZN(n2165) );
  XNOR2_X2 U4225 ( .A(n2169), .B(n2714), .ZN(n2279) );
  NAND2_X2 U4226 ( .A1(n2967), .A2(n3223), .ZN(n2169) );
  NAND2_X1 U4227 ( .A1(n1524), .A2(n3840), .ZN(n3841) );
  NAND2_X1 U4228 ( .A1(n1524), .A2(n2706), .ZN(n3649) );
  NAND2_X1 U4229 ( .A1(n1524), .A2(n4317), .ZN(n4318) );
  NAND2_X1 U4230 ( .A1(n1524), .A2(n3796), .ZN(n3798) );
  NAND2_X1 U4231 ( .A1(n1524), .A2(n3785), .ZN(n3786) );
  INV_X2 U4232 ( .A(n4249), .ZN(n3035) );
  NAND2_X2 U4233 ( .A1(b[0]), .A2(n1326), .ZN(n4249) );
  NAND2_X2 U4234 ( .A1(n2490), .A2(n965), .ZN(n2170) );
  INV_X4 U4235 ( .A(n2427), .ZN(n4280) );
  AOI22_X2 U4236 ( .A1(n4570), .A2(n6293), .B1(n4565), .B2(n4569), .ZN(n4571)
         );
  NAND2_X4 U4237 ( .A1(n2271), .A2(n2270), .ZN(n4564) );
  NOR2_X2 U4238 ( .A1(n3051), .A2(n1004), .ZN(n2181) );
  INV_X2 U4239 ( .A(n4484), .ZN(n2182) );
  INV_X4 U4240 ( .A(n4464), .ZN(n2184) );
  NAND2_X2 U4241 ( .A1(n2186), .A2(n2185), .ZN(n4213) );
  NOR2_X2 U4242 ( .A1(n4236), .A2(n6569), .ZN(n2187) );
  INV_X4 U4243 ( .A(n3227), .ZN(n2194) );
  NOR2_X2 U4244 ( .A1(n2748), .A2(n3888), .ZN(n2195) );
  XNOR2_X2 U4246 ( .A(n5238), .B(n5290), .ZN(n5307) );
  NAND3_X2 U4247 ( .A1(n1659), .A2(n3115), .A3(n987), .ZN(n2200) );
  NOR2_X1 U4251 ( .A1(n4774), .A2(n5105), .ZN(n2203) );
  NOR2_X2 U4252 ( .A1(n3161), .A2(b[22]), .ZN(n2204) );
  NAND2_X2 U4253 ( .A1(n2207), .A2(n2206), .ZN(n2205) );
  NAND2_X2 U4255 ( .A1(n3697), .A2(n5247), .ZN(n2207) );
  NAND2_X2 U4256 ( .A1(n3423), .A2(n958), .ZN(n4279) );
  NAND2_X2 U4257 ( .A1(n3301), .A2(n3857), .ZN(n2209) );
  NAND2_X2 U4259 ( .A1(n2214), .A2(n2211), .ZN(n3859) );
  NAND2_X2 U4261 ( .A1(n3821), .A2(n3822), .ZN(n2214) );
  INV_X8 U4263 ( .A(a[5]), .ZN(n4821) );
  NAND2_X2 U4264 ( .A1(n2217), .A2(n2216), .ZN(n3291) );
  NAND2_X2 U4266 ( .A1(n3293), .A2(n3292), .ZN(n2217) );
  OAI21_X2 U4268 ( .B1(n5079), .B2(n4359), .A(n6455), .ZN(n4444) );
  NAND2_X2 U4271 ( .A1(n4033), .A2(n6191), .ZN(n2223) );
  NOR2_X2 U4273 ( .A1(n2543), .A2(n1057), .ZN(n2224) );
  NAND2_X1 U4274 ( .A1(n3865), .A2(n6459), .ZN(n2225) );
  OAI21_X2 U4275 ( .B1(n1003), .B2(n751), .A(n3082), .ZN(n4635) );
  NAND2_X2 U4276 ( .A1(n2228), .A2(n2227), .ZN(n2229) );
  INV_X2 U4277 ( .A(n3446), .ZN(n2227) );
  NAND2_X2 U4278 ( .A1(n2375), .A2(n6366), .ZN(n2228) );
  INV_X2 U4280 ( .A(n2956), .ZN(n2232) );
  NAND2_X2 U4282 ( .A1(n5647), .A2(n4148), .ZN(n5657) );
  XNOR2_X2 U4283 ( .A(n2233), .B(n4139), .ZN(n5647) );
  XNOR2_X2 U4284 ( .A(n4141), .B(n4142), .ZN(n2233) );
  NAND2_X2 U4285 ( .A1(n2234), .A2(n5648), .ZN(n4148) );
  NAND2_X2 U4286 ( .A1(n5649), .A2(n5650), .ZN(n2234) );
  NAND3_X2 U4287 ( .A1(n3274), .A2(n2236), .A3(n2293), .ZN(n3732) );
  NAND2_X2 U4288 ( .A1(n1021), .A2(n2235), .ZN(n2293) );
  INV_X2 U4290 ( .A(n3534), .ZN(n2237) );
  NAND2_X4 U4293 ( .A1(n2295), .A2(n3275), .ZN(n5733) );
  NAND2_X2 U4294 ( .A1(n2241), .A2(n4305), .ZN(n3212) );
  NAND2_X2 U4295 ( .A1(n2240), .A2(n4276), .ZN(n2239) );
  INV_X2 U4296 ( .A(n4274), .ZN(n2240) );
  INV_X2 U4298 ( .A(n3356), .ZN(n2242) );
  NAND2_X2 U4299 ( .A1(n2450), .A2(n4765), .ZN(n2449) );
  BUF_X4 U4300 ( .A(n4765), .Z(n2243) );
  NAND2_X2 U4302 ( .A1(n782), .A2(n4181), .ZN(n4229) );
  NAND2_X2 U4303 ( .A1(n2246), .A2(n2245), .ZN(n4180) );
  NAND2_X2 U4304 ( .A1(n3358), .A2(b[3]), .ZN(n2245) );
  NOR2_X2 U4306 ( .A1(n4800), .A2(b[3]), .ZN(n2250) );
  NOR2_X2 U4307 ( .A1(n2253), .A2(n2252), .ZN(n2251) );
  NAND2_X2 U4310 ( .A1(n2260), .A2(n2259), .ZN(n2258) );
  OAI21_X2 U4311 ( .B1(n3867), .B2(n3868), .A(n3912), .ZN(n2259) );
  NAND2_X2 U4312 ( .A1(n3183), .A2(n460), .ZN(n2260) );
  NOR2_X2 U4313 ( .A1(n3186), .A2(n3910), .ZN(n2263) );
  INV_X2 U4314 ( .A(n4119), .ZN(n4120) );
  NAND2_X2 U4315 ( .A1(n2264), .A2(b[0]), .ZN(n4119) );
  INV_X1 U4316 ( .A(n505), .ZN(n2264) );
  NOR2_X1 U4317 ( .A1(n5746), .A2(n2265), .ZN(n5741) );
  AOI21_X1 U4318 ( .B1(n5728), .B2(n2265), .A(n5746), .ZN(n5732) );
  NAND2_X1 U4320 ( .A1(n5783), .A2(n710), .ZN(n5784) );
  OAI21_X1 U4321 ( .B1(n5797), .B2(n5796), .A(n710), .ZN(n5802) );
  INV_X2 U4322 ( .A(n3316), .ZN(n2268) );
  NOR2_X4 U4323 ( .A1(n2269), .A2(n5598), .ZN(n5968) );
  NAND2_X4 U4324 ( .A1(n2269), .A2(n5598), .ZN(n5599) );
  XNOR2_X1 U4325 ( .A(n5598), .B(n2269), .ZN(n2705) );
  NAND2_X4 U4326 ( .A1(n3471), .A2(n3498), .ZN(n2269) );
  INV_X2 U4330 ( .A(n3899), .ZN(n2277) );
  AOI21_X2 U4332 ( .B1(n5380), .B2(n2278), .A(n5379), .ZN(n5625) );
  NAND2_X2 U4333 ( .A1(n5381), .A2(n2278), .ZN(n5382) );
  NOR2_X2 U4334 ( .A1(n3380), .A2(n3714), .ZN(n2282) );
  NAND2_X2 U4335 ( .A1(n2777), .A2(n3381), .ZN(n3714) );
  NAND2_X4 U4336 ( .A1(n2284), .A2(a[15]), .ZN(n5219) );
  NOR2_X2 U4337 ( .A1(n3848), .A2(n2288), .ZN(n2287) );
  NOR2_X2 U4338 ( .A1(n4810), .A2(n1324), .ZN(n2288) );
  OAI21_X2 U4344 ( .B1(n1107), .B2(n3540), .A(n5422), .ZN(n2587) );
  INV_X2 U4346 ( .A(n3200), .ZN(n2317) );
  NAND2_X2 U4349 ( .A1(n2862), .A2(n6133), .ZN(n6131) );
  INV_X2 U4351 ( .A(n5938), .ZN(n2332) );
  XNOR2_X2 U4352 ( .A(n2437), .B(n3887), .ZN(n2334) );
  NOR2_X4 U4355 ( .A1(n2338), .A2(n5372), .ZN(n5571) );
  NAND2_X2 U4356 ( .A1(n4158), .A2(n4157), .ZN(n4194) );
  NAND2_X2 U4357 ( .A1(n2341), .A2(n2340), .ZN(n5563) );
  NAND3_X1 U4358 ( .A1(n966), .A2(n5550), .A3(n2344), .ZN(n2340) );
  INV_X2 U4359 ( .A(n2342), .ZN(n2341) );
  AOI21_X2 U4360 ( .B1(n966), .B2(n2344), .A(n5550), .ZN(n2342) );
  XNOR2_X2 U4361 ( .A(n5497), .B(n5496), .ZN(n2345) );
  NOR2_X2 U4362 ( .A1(n2343), .A2(n5346), .ZN(n5492) );
  INV_X2 U4363 ( .A(n5348), .ZN(n2343) );
  INV_X2 U4364 ( .A(n2344), .ZN(n5549) );
  NAND2_X2 U4365 ( .A1(n2345), .A2(n5501), .ZN(n2344) );
  AOI21_X2 U4366 ( .B1(n3508), .B2(n265), .A(n2347), .ZN(n2346) );
  INV_X2 U4368 ( .A(n2354), .ZN(n2352) );
  NAND3_X2 U4370 ( .A1(n3451), .A2(n5113), .A3(n3450), .ZN(n2360) );
  NAND2_X2 U4371 ( .A1(n2359), .A2(n2357), .ZN(n2356) );
  INV_X2 U4372 ( .A(n5080), .ZN(n2358) );
  INV_X2 U4373 ( .A(n2489), .ZN(n2359) );
  INV_X2 U4374 ( .A(n5081), .ZN(n2361) );
  OAI21_X2 U4375 ( .B1(n5083), .B2(n5081), .A(n5082), .ZN(n2362) );
  NOR2_X1 U4376 ( .A1(n5081), .A2(n3690), .ZN(n2363) );
  AOI21_X1 U4377 ( .B1(n5711), .B2(n6180), .A(n5710), .ZN(n5715) );
  NAND2_X2 U4378 ( .A1(n3042), .A2(n3041), .ZN(n4470) );
  AOI21_X2 U4379 ( .B1(n4820), .B2(n1287), .A(n4819), .ZN(n4872) );
  AOI22_X2 U4380 ( .A1(n3066), .A2(n4873), .B1(n2370), .B2(n3556), .ZN(n2369)
         );
  INV_X4 U4384 ( .A(n3341), .ZN(n5092) );
  NOR2_X2 U4386 ( .A1(n4191), .A2(n4190), .ZN(n2377) );
  NAND3_X2 U4387 ( .A1(n4045), .A2(a[9]), .A3(n4998), .ZN(n4999) );
  INV_X2 U4388 ( .A(n2379), .ZN(n2378) );
  NAND2_X2 U4389 ( .A1(n4544), .A2(a[9]), .ZN(n2379) );
  NAND2_X2 U4390 ( .A1(n5182), .A2(n2953), .ZN(n3697) );
  NAND2_X2 U4391 ( .A1(n5178), .A2(n3562), .ZN(n2953) );
  INV_X8 U4392 ( .A(n3673), .ZN(n3562) );
  AOI21_X2 U4393 ( .B1(n2380), .B2(n5266), .A(n5181), .ZN(n5182) );
  INV_X2 U4394 ( .A(n2381), .ZN(n3553) );
  NAND3_X2 U4395 ( .A1(n3770), .A2(n4987), .A3(n2381), .ZN(n5098) );
  NAND2_X2 U4396 ( .A1(n2382), .A2(b[10]), .ZN(n3295) );
  NAND2_X2 U4397 ( .A1(n2382), .A2(b[0]), .ZN(n3908) );
  MUX2_X2 U4399 ( .A(n2382), .B(n2510), .S(n5951), .Z(n5341) );
  INV_X8 U4401 ( .A(n5423), .ZN(n2382) );
  NAND3_X1 U4402 ( .A1(n2384), .A2(n1844), .A3(n2488), .ZN(n2461) );
  NAND2_X2 U4403 ( .A1(n3119), .A2(n991), .ZN(n4078) );
  NAND3_X2 U4405 ( .A1(n2387), .A2(n3119), .A3(n991), .ZN(n2385) );
  INV_X2 U4406 ( .A(n4008), .ZN(n2387) );
  NAND2_X2 U4407 ( .A1(n2390), .A2(n2388), .ZN(n3398) );
  INV_X2 U4408 ( .A(n2575), .ZN(n2390) );
  NAND2_X2 U4411 ( .A1(n2395), .A2(n2394), .ZN(n4842) );
  NAND2_X2 U4412 ( .A1(n5947), .A2(n1324), .ZN(n2394) );
  NAND2_X2 U4413 ( .A1(n5900), .A2(b[6]), .ZN(n2395) );
  INV_X2 U4414 ( .A(n5063), .ZN(n5066) );
  NAND2_X2 U4415 ( .A1(n2397), .A2(n2396), .ZN(n5063) );
  NAND2_X2 U4416 ( .A1(n5024), .A2(n985), .ZN(n2396) );
  INV_X2 U4417 ( .A(n2398), .ZN(n5319) );
  NOR2_X2 U4418 ( .A1(n2400), .A2(n3413), .ZN(n2399) );
  INV_X2 U4420 ( .A(n3598), .ZN(n3334) );
  INV_X2 U4421 ( .A(n4338), .ZN(n3580) );
  XNOR2_X2 U4423 ( .A(n5226), .B(n5229), .ZN(n2404) );
  BUF_X4 U4425 ( .A(n5423), .Z(n2406) );
  NAND2_X2 U4426 ( .A1(n2408), .A2(n2407), .ZN(n5119) );
  AOI22_X2 U4427 ( .A1(n309), .A2(b[17]), .B1(b[16]), .B2(n2406), .ZN(n2407)
         );
  NOR2_X4 U4428 ( .A1(n3688), .A2(n3686), .ZN(n2826) );
  AOI22_X2 U4429 ( .A1(n2666), .A2(n2667), .B1(n4631), .B2(n4632), .ZN(n2411)
         );
  NAND3_X2 U4431 ( .A1(n790), .A2(n6303), .A3(n3382), .ZN(n2414) );
  NAND3_X2 U4433 ( .A1(n2420), .A2(n2426), .A3(n3350), .ZN(n2419) );
  NAND2_X2 U4438 ( .A1(n3376), .A2(n5037), .ZN(n2425) );
  INV_X2 U4439 ( .A(n4270), .ZN(n2430) );
  OAI22_X2 U4440 ( .A1(n606), .A2(n2249), .B1(n513), .B2(b[2]), .ZN(n2431) );
  NOR2_X2 U4441 ( .A1(n2433), .A2(n3598), .ZN(n2593) );
  XNOR2_X2 U4442 ( .A(b[11]), .B(a[21]), .ZN(n2433) );
  NAND2_X4 U4447 ( .A1(n2455), .A2(n2454), .ZN(n3304) );
  NAND2_X2 U4448 ( .A1(n608), .A2(n6529), .ZN(n2454) );
  OAI21_X2 U4449 ( .B1(n2460), .B2(n2467), .A(n2459), .ZN(n2456) );
  INV_X2 U4451 ( .A(n4620), .ZN(n2462) );
  NAND2_X4 U4456 ( .A1(n2473), .A2(a[13]), .ZN(n4940) );
  OAI21_X2 U4457 ( .B1(n2281), .B2(n3380), .A(n2475), .ZN(n2998) );
  INV_X2 U4458 ( .A(n3714), .ZN(n2475) );
  NAND2_X2 U4459 ( .A1(n2477), .A2(n2476), .ZN(n5086) );
  NAND2_X2 U4460 ( .A1(n5028), .A2(n5027), .ZN(n2476) );
  NAND3_X2 U4464 ( .A1(n6151), .A2(n2491), .A3(n3491), .ZN(n2482) );
  NAND2_X2 U4468 ( .A1(n2955), .A2(n2493), .ZN(n3360) );
  NAND2_X1 U4469 ( .A1(n5972), .A2(n2493), .ZN(n5977) );
  NAND2_X2 U4470 ( .A1(n5318), .A2(n5319), .ZN(n2493) );
  NAND2_X2 U4471 ( .A1(n2494), .A2(n2495), .ZN(n5308) );
  OAI21_X1 U4472 ( .B1(n2499), .B2(n5263), .A(n2497), .ZN(n2494) );
  NAND2_X2 U4473 ( .A1(n5265), .A2(n2496), .ZN(n2495) );
  NOR2_X1 U4474 ( .A1(n5263), .A2(n2497), .ZN(n2496) );
  NAND2_X2 U4476 ( .A1(n2502), .A2(n2501), .ZN(n2500) );
  NAND3_X2 U4477 ( .A1(n2504), .A2(n2982), .A3(n3611), .ZN(\d[41]_BAR ) );
  INV_X2 U4478 ( .A(n2505), .ZN(n2504) );
  NAND2_X2 U4479 ( .A1(n6012), .A2(n2981), .ZN(n2505) );
  INV_X8 U4482 ( .A(n4768), .ZN(n2510) );
  NAND2_X2 U4483 ( .A1(n5058), .A2(n5057), .ZN(n2512) );
  BUF_X4 U4484 ( .A(n4829), .Z(n2514) );
  MUX2_X2 U4485 ( .A(n2514), .B(n5526), .S(n5951), .Z(n5411) );
  MUX2_X2 U4486 ( .A(n2514), .B(n5526), .S(n5360), .Z(n5440) );
  NAND2_X2 U4487 ( .A1(n2515), .A2(n5727), .ZN(n2638) );
  NOR2_X2 U4488 ( .A1(n5060), .A2(n5061), .ZN(n2517) );
  AOI21_X2 U4490 ( .B1(n5556), .B2(n5557), .A(n5555), .ZN(n5561) );
  NOR2_X2 U4491 ( .A1(n2522), .A2(n2520), .ZN(n5555) );
  AOI22_X2 U4492 ( .A1(n2521), .A2(n5370), .B1(n6508), .B2(n5368), .ZN(n2520)
         );
  NAND2_X2 U4493 ( .A1(n2812), .A2(n5367), .ZN(n2521) );
  NAND2_X1 U4497 ( .A1(n4829), .A2(b[6]), .ZN(n2525) );
  NAND2_X2 U4498 ( .A1(n4742), .A2(n585), .ZN(n2527) );
  NAND2_X2 U4499 ( .A1(n4583), .A2(n2529), .ZN(n5823) );
  NAND2_X2 U4500 ( .A1(n3978), .A2(n3977), .ZN(n4075) );
  MUX2_X2 U4506 ( .A(n5409), .B(n2537), .S(b[23]), .Z(n5410) );
  MUX2_X2 U4507 ( .A(n2537), .B(n5266), .S(n5529), .Z(n5269) );
  MUX2_X2 U4509 ( .A(n2537), .B(n6524), .S(n981), .Z(n4898) );
  MUX2_X2 U4510 ( .A(n2537), .B(n5266), .S(n5951), .Z(n5426) );
  MUX2_X2 U4511 ( .A(n2537), .B(n6524), .S(n5105), .Z(n5396) );
  MUX2_X2 U4512 ( .A(n2537), .B(n6524), .S(n5471), .Z(n5467) );
  INV_X8 U4513 ( .A(n5179), .ZN(n2537) );
  INV_X4 U4515 ( .A(n4636), .ZN(n2539) );
  INV_X2 U4519 ( .A(n3357), .ZN(n2553) );
  NAND2_X2 U4520 ( .A1(n2557), .A2(n2554), .ZN(n5280) );
  NAND3_X2 U4521 ( .A1(n2558), .A2(n2557), .A3(n2554), .ZN(n5356) );
  NAND2_X2 U4522 ( .A1(n3661), .A2(n2555), .ZN(n2554) );
  INV_X2 U4523 ( .A(n2556), .ZN(n2555) );
  NAND2_X2 U4524 ( .A1(n5351), .A2(n5349), .ZN(n2556) );
  NAND2_X2 U4526 ( .A1(n2560), .A2(n2559), .ZN(n5281) );
  INV_X2 U4527 ( .A(n2561), .ZN(n2560) );
  INV_X2 U4528 ( .A(n5279), .ZN(n2562) );
  NAND2_X4 U4529 ( .A1(n2563), .A2(a[1]), .ZN(n4491) );
  INV_X8 U4530 ( .A(a[0]), .ZN(n2563) );
  NAND2_X2 U4531 ( .A1(n2566), .A2(n6239), .ZN(n2565) );
  INV_X2 U4533 ( .A(n3093), .ZN(n2677) );
  NAND2_X2 U4534 ( .A1(n2674), .A2(n2673), .ZN(n2573) );
  NAND2_X4 U4536 ( .A1(n366), .A2(n5316), .ZN(n5597) );
  NAND3_X2 U4537 ( .A1(n2575), .A2(n3588), .A3(n3589), .ZN(n3397) );
  INV_X1 U4538 ( .A(n4415), .ZN(n5337) );
  XNOR2_X2 U4541 ( .A(n1417), .B(n2758), .ZN(n2582) );
  INV_X4 U4542 ( .A(n2583), .ZN(n4634) );
  NAND2_X2 U4543 ( .A1(n3398), .A2(n3397), .ZN(n2583) );
  NOR2_X2 U4544 ( .A1(n3104), .A2(n4924), .ZN(n2584) );
  OAI22_X2 U4545 ( .A1(n606), .A2(n5951), .B1(n512), .B2(b[21]), .ZN(n2585) );
  NAND2_X2 U4546 ( .A1(n5573), .A2(n5572), .ZN(n5995) );
  NAND2_X4 U4547 ( .A1(a[17]), .A2(a[18]), .ZN(n2954) );
  AOI22_X2 U4549 ( .A1(n1761), .A2(n4942), .B1(n5136), .B2(b[10]), .ZN(n2594)
         );
  INV_X4 U4550 ( .A(n2597), .ZN(n2600) );
  NAND2_X2 U4551 ( .A1(n3092), .A2(n3091), .ZN(n5034) );
  NAND2_X2 U4552 ( .A1(n3091), .A2(n3092), .ZN(n2598) );
  NAND2_X2 U4554 ( .A1(n2605), .A2(n2606), .ZN(n2604) );
  OAI21_X2 U4556 ( .B1(n2611), .B2(n4580), .A(n2610), .ZN(n2609) );
  NOR2_X2 U4558 ( .A1(n2616), .A2(n4517), .ZN(n2615) );
  NAND2_X2 U4559 ( .A1(n2618), .A2(n2617), .ZN(n2616) );
  NAND3_X2 U4562 ( .A1(n2620), .A2(n4512), .A3(n4515), .ZN(n2619) );
  NAND2_X2 U4563 ( .A1(n4516), .A2(n4514), .ZN(n2620) );
  NAND2_X4 U4566 ( .A1(n2912), .A2(n2911), .ZN(n3673) );
  XNOR2_X2 U4567 ( .A(b[7]), .B(a[19]), .ZN(n2621) );
  NAND2_X2 U4570 ( .A1(n2625), .A2(n2624), .ZN(n4968) );
  NAND2_X2 U4571 ( .A1(n3315), .A2(n2626), .ZN(n2625) );
  NAND2_X2 U4572 ( .A1(n2627), .A2(n2628), .ZN(n2626) );
  NOR2_X4 U4573 ( .A1(n3252), .A2(n4884), .ZN(n2629) );
  OAI22_X2 U4574 ( .A1(n5477), .A2(b[3]), .B1(n3538), .B2(n4752), .ZN(n2632)
         );
  NOR2_X2 U4576 ( .A1(n4866), .A2(n4865), .ZN(n2634) );
  NAND2_X2 U4577 ( .A1(n3316), .A2(n4638), .ZN(n2899) );
  NAND3_X2 U4578 ( .A1(n5772), .A2(n2742), .A3(n4316), .ZN(n5727) );
  NAND2_X2 U4581 ( .A1(a[5]), .A2(n979), .ZN(n2642) );
  NAND2_X2 U4582 ( .A1(n4821), .A2(b[23]), .ZN(n2643) );
  AOI21_X2 U4586 ( .B1(n4345), .B2(n4447), .A(n2648), .ZN(n4374) );
  BUF_X4 U4587 ( .A(n452), .Z(n2650) );
  NOR2_X2 U4588 ( .A1(n3042), .A2(n3041), .ZN(n3347) );
  NAND2_X1 U4592 ( .A1(n5086), .A2(n5087), .ZN(n2655) );
  INV_X8 U4593 ( .A(n5076), .ZN(n2656) );
  NAND2_X1 U4597 ( .A1(n5284), .A2(n5283), .ZN(n2660) );
  INV_X2 U4600 ( .A(n3517), .ZN(n2662) );
  NAND2_X1 U4601 ( .A1(n2861), .A2(n5565), .ZN(n2665) );
  NOR2_X1 U4605 ( .A1(b[15]), .A2(n568), .ZN(n3963) );
  NAND2_X4 U4606 ( .A1(n3633), .A2(n4999), .ZN(n5042) );
  NAND2_X1 U4608 ( .A1(n3986), .A2(n3985), .ZN(n2668) );
  NAND2_X1 U4609 ( .A1(n3823), .A2(n3813), .ZN(n2670) );
  NAND2_X1 U4610 ( .A1(n3814), .A2(n3813), .ZN(n2671) );
  NAND2_X1 U4611 ( .A1(n3814), .A2(n3823), .ZN(n2672) );
  NAND3_X2 U4612 ( .A1(n2672), .A2(n2671), .A3(n2670), .ZN(n3861) );
  NOR2_X1 U4615 ( .A1(n3492), .A2(n4581), .ZN(n4644) );
  INV_X1 U4616 ( .A(n5034), .ZN(n5031) );
  INV_X4 U4618 ( .A(n628), .ZN(n3689) );
  INV_X2 U4619 ( .A(n3150), .ZN(n2678) );
  INV_X1 U4620 ( .A(n4803), .ZN(n2679) );
  NAND2_X1 U4621 ( .A1(n5629), .A2(n637), .ZN(n5975) );
  INV_X1 U4622 ( .A(n565), .ZN(n2680) );
  NAND2_X4 U4623 ( .A1(a[12]), .A2(a[11]), .ZN(n2686) );
  NAND2_X4 U4624 ( .A1(n2684), .A2(n2685), .ZN(n2687) );
  NAND2_X4 U4625 ( .A1(n2687), .A2(n2686), .ZN(n4010) );
  INV_X8 U4627 ( .A(a[11]), .ZN(n2685) );
  NAND2_X4 U4629 ( .A1(a[1]), .A2(a[2]), .ZN(n2697) );
  NAND2_X4 U4630 ( .A1(n2695), .A2(n2696), .ZN(n2698) );
  NAND2_X4 U4631 ( .A1(n2698), .A2(n2697), .ZN(n3484) );
  INV_X8 U4632 ( .A(a[1]), .ZN(n2695) );
  INV_X8 U4633 ( .A(a[2]), .ZN(n2696) );
  NAND2_X1 U4634 ( .A1(n4494), .A2(n6215), .ZN(n3187) );
  INV_X8 U4635 ( .A(b[10]), .ZN(n4942) );
  INV_X8 U4636 ( .A(a[20]), .ZN(n2699) );
  OR2_X4 U4637 ( .A1(n3597), .A2(n3598), .ZN(n3599) );
  NAND2_X1 U4638 ( .A1(n3367), .A2(n5473), .ZN(n3243) );
  OAI21_X1 U4639 ( .B1(n3326), .B2(n5104), .A(n5166), .ZN(n3027) );
  AOI21_X1 U4640 ( .B1(n5076), .B2(n5951), .A(n3505), .ZN(n3504) );
  NAND2_X1 U4641 ( .A1(n953), .A2(n5221), .ZN(n5222) );
  OAI21_X1 U4642 ( .B1(n4250), .B2(n4249), .A(n3320), .ZN(n4252) );
  NAND2_X1 U4643 ( .A1(n6040), .A2(n3154), .ZN(n6034) );
  BUF_X4 U4645 ( .A(n2899), .Z(n2988) );
  INV_X1 U4646 ( .A(n6124), .ZN(n6120) );
  NOR2_X1 U4647 ( .A1(n4309), .A2(n4308), .ZN(n4310) );
  INV_X1 U4648 ( .A(n5823), .ZN(n5814) );
  NAND2_X1 U4649 ( .A1(n5824), .A2(n6453), .ZN(n5827) );
  INV_X1 U4650 ( .A(n6206), .ZN(n3098) );
  OAI21_X1 U4653 ( .B1(n1358), .B2(n4678), .A(n4673), .ZN(n4676) );
  INV_X1 U4654 ( .A(n4724), .ZN(n4673) );
  NOR2_X1 U4655 ( .A1(n5104), .A2(n5166), .ZN(n3472) );
  NOR2_X1 U4656 ( .A1(n5952), .A2(b[5]), .ZN(n4843) );
  NOR2_X1 U4657 ( .A1(n6457), .A2(b[11]), .ZN(n3652) );
  INV_X1 U4660 ( .A(n4761), .ZN(n3128) );
  NAND2_X2 U4663 ( .A1(n5951), .A2(a[3]), .ZN(n4697) );
  NOR2_X1 U4664 ( .A1(n5110), .A2(n5293), .ZN(n4756) );
  NOR2_X1 U4665 ( .A1(n3572), .A2(n5218), .ZN(n3413) );
  NOR2_X1 U4666 ( .A1(n4829), .A2(n2143), .ZN(n4832) );
  INV_X1 U4668 ( .A(n5104), .ZN(n3241) );
  NOR2_X1 U4669 ( .A1(n3445), .A2(n1896), .ZN(n2915) );
  NAND2_X1 U4670 ( .A1(n5422), .A2(n1896), .ZN(n3490) );
  NOR2_X1 U4671 ( .A1(n5445), .A2(b[0]), .ZN(n3781) );
  NAND2_X1 U4672 ( .A1(n6155), .A2(n984), .ZN(n3566) );
  INV_X1 U4673 ( .A(n4448), .ZN(n4440) );
  INV_X1 U4674 ( .A(n5123), .ZN(n5121) );
  INV_X1 U4676 ( .A(n5062), .ZN(n5067) );
  NOR2_X1 U4677 ( .A1(n5063), .A2(n5064), .ZN(n5068) );
  NAND2_X1 U4678 ( .A1(n3445), .A2(b[18]), .ZN(n3309) );
  NAND2_X1 U4679 ( .A1(n3351), .A2(n3438), .ZN(n2819) );
  NAND2_X1 U4680 ( .A1(n47), .A2(b[0]), .ZN(n3702) );
  NAND3_X1 U4681 ( .A1(n4948), .A2(a[7]), .A3(n248), .ZN(n4082) );
  NAND3_X1 U4684 ( .A1(n4204), .A2(n6178), .A3(n4205), .ZN(n4206) );
  INV_X1 U4685 ( .A(n5670), .ZN(n4204) );
  INV_X1 U4686 ( .A(n4383), .ZN(n4386) );
  NOR2_X1 U4691 ( .A1(n5498), .A2(n5952), .ZN(n5499) );
  AOI22_X1 U4692 ( .A1(n5317), .A2(n5309), .B1(n1001), .B2(n5308), .ZN(n5318)
         );
  INV_X1 U4694 ( .A(n4101), .ZN(n4096) );
  NAND2_X1 U4695 ( .A1(n4070), .A2(n818), .ZN(n2972) );
  INV_X1 U4696 ( .A(n4644), .ZN(n4645) );
  NAND2_X1 U4700 ( .A1(n5958), .A2(n5957), .ZN(n5960) );
  INV_X1 U4701 ( .A(n6121), .ZN(n6123) );
  INV_X1 U4702 ( .A(n6122), .ZN(n6119) );
  NOR2_X1 U4703 ( .A1(n6104), .A2(n5952), .ZN(n6105) );
  INV_X1 U4704 ( .A(n4260), .ZN(n4263) );
  NAND2_X1 U4705 ( .A1(n4260), .A2(n6201), .ZN(n4264) );
  NAND2_X1 U4707 ( .A1(n4635), .A2(n4636), .ZN(n3447) );
  AOI21_X1 U4708 ( .B1(n6376), .B2(n2938), .A(n2937), .ZN(n3005) );
  NAND2_X1 U4710 ( .A1(n5379), .A2(n2782), .ZN(n2780) );
  INV_X1 U4711 ( .A(n5981), .ZN(n5982) );
  INV_X1 U4713 ( .A(n6063), .ZN(n5576) );
  NAND2_X1 U4714 ( .A1(n6075), .A2(n6065), .ZN(n6066) );
  INV_X1 U4715 ( .A(n6064), .ZN(n6067) );
  NAND2_X1 U4716 ( .A1(n6112), .A2(n6117), .ZN(n6108) );
  NAND3_X1 U4717 ( .A1(n472), .A2(n4125), .A3(n3540), .ZN(n4127) );
  XNOR2_X1 U4718 ( .A(n6097), .B(n6096), .ZN(n6099) );
  NAND2_X1 U4719 ( .A1(n5648), .A2(n5649), .ZN(n6098) );
  INV_X1 U4720 ( .A(n5650), .ZN(n5651) );
  XNOR2_X1 U4721 ( .A(n163), .B(n5648), .ZN(n5654) );
  NAND2_X1 U4722 ( .A1(n5656), .A2(n5657), .ZN(n5659) );
  INV_X1 U4723 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U4725 ( .A1(n4117), .A2(n4116), .ZN(n4112) );
  NOR2_X1 U4727 ( .A1(n5693), .A2(n5689), .ZN(n4234) );
  NAND2_X1 U4728 ( .A1(n5693), .A2(n5689), .ZN(n4233) );
  NOR2_X1 U4729 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  NAND2_X1 U4730 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  NAND2_X1 U4731 ( .A1(n5773), .A2(n5772), .ZN(n5775) );
  NOR3_X1 U4732 ( .A1(n5750), .A2(n5778), .A3(n5747), .ZN(n5744) );
  OAI22_X1 U4733 ( .A1(n5747), .A2(n6522), .B1(n5783), .B2(n5748), .ZN(n5743)
         );
  INV_X1 U4734 ( .A(n5747), .ZN(n5751) );
  NAND3_X1 U4735 ( .A1(n5758), .A2(n5753), .A3(n5778), .ZN(n5754) );
  XNOR2_X1 U4737 ( .A(n976), .B(n5799), .ZN(n5800) );
  NOR2_X1 U4738 ( .A1(n5792), .A2(n5791), .ZN(n5803) );
  INV_X1 U4740 ( .A(n5837), .ZN(n5849) );
  INV_X1 U4743 ( .A(n5605), .ZN(n5606) );
  NAND3_X1 U4744 ( .A1(n6025), .A2(n5963), .A3(n2851), .ZN(n5966) );
  INV_X1 U4745 ( .A(n5964), .ZN(n5963) );
  NAND2_X1 U4746 ( .A1(n5952), .A2(b[6]), .ZN(n4813) );
  NAND2_X1 U4747 ( .A1(n3639), .A2(b[9]), .ZN(n3959) );
  INV_X1 U4748 ( .A(n4948), .ZN(n3878) );
  NAND2_X1 U4752 ( .A1(n3058), .A2(b[12]), .ZN(n3056) );
  NAND2_X1 U4753 ( .A1(n2730), .A2(n1059), .ZN(n3071) );
  NOR2_X1 U4754 ( .A1(n4504), .A2(n3438), .ZN(n3437) );
  NOR2_X1 U4756 ( .A1(n4834), .A2(b[23]), .ZN(n4675) );
  NAND2_X1 U4757 ( .A1(n3470), .A2(n4729), .ZN(n3246) );
  NAND2_X1 U4758 ( .A1(n5277), .A2(n5266), .ZN(n4944) );
  NOR2_X1 U4761 ( .A1(n4601), .A2(n981), .ZN(n3653) );
  NOR2_X1 U4762 ( .A1(n3969), .A2(n4490), .ZN(n3343) );
  NOR2_X1 U4763 ( .A1(n5077), .A2(n4598), .ZN(n4053) );
  NOR2_X1 U4764 ( .A1(n3617), .A2(n3054), .ZN(n3053) );
  NAND2_X1 U4765 ( .A1(n3058), .A2(b[11]), .ZN(n3054) );
  INV_X1 U4767 ( .A(n4061), .ZN(n4062) );
  NOR2_X1 U4769 ( .A1(n3540), .A2(n3598), .ZN(n4429) );
  NOR2_X1 U4772 ( .A1(n760), .A2(n1324), .ZN(n4498) );
  NOR2_X1 U4774 ( .A1(n465), .A2(n3342), .ZN(n2836) );
  NOR2_X2 U4776 ( .A1(n3699), .A2(n4825), .ZN(n4827) );
  NAND2_X1 U4777 ( .A1(n5525), .A2(b[19]), .ZN(n2820) );
  NOR2_X1 U4779 ( .A1(n3699), .A2(n3442), .ZN(n3441) );
  NAND2_X1 U4780 ( .A1(a[19]), .A2(n5105), .ZN(n3442) );
  AOI21_X1 U4781 ( .B1(n3263), .B2(n2380), .A(n5952), .ZN(n5398) );
  NOR2_X1 U4783 ( .A1(n805), .A2(n3367), .ZN(n3543) );
  NOR2_X1 U4784 ( .A1(n3538), .A2(n4590), .ZN(n3776) );
  NOR2_X1 U4785 ( .A1(n6211), .A2(n984), .ZN(n3964) );
  NAND2_X1 U4786 ( .A1(n3975), .A2(n3976), .ZN(n2866) );
  OAI21_X1 U4787 ( .B1(n3976), .B2(n3975), .A(n3974), .ZN(n2867) );
  NAND2_X1 U4788 ( .A1(n4453), .A2(n2919), .ZN(n4454) );
  NOR2_X1 U4790 ( .A1(b[2]), .A2(n5473), .ZN(n3177) );
  AOI22_X1 U4791 ( .A1(n4810), .A2(b[14]), .B1(n5293), .B2(n4746), .ZN(n3577)
         );
  NAND2_X1 U4792 ( .A1(n4021), .A2(n5471), .ZN(n4494) );
  NAND2_X1 U4795 ( .A1(n4616), .A2(n4617), .ZN(n4620) );
  INV_X1 U4797 ( .A(n5052), .ZN(n5055) );
  NAND2_X1 U4799 ( .A1(n5246), .A2(n5247), .ZN(n5249) );
  NAND2_X1 U4800 ( .A1(n5277), .A2(a[23]), .ZN(n5278) );
  INV_X1 U4801 ( .A(n5445), .ZN(n5442) );
  NOR2_X1 U4802 ( .A1(n3699), .A2(n4896), .ZN(n4897) );
  NAND3_X1 U4804 ( .A1(n3488), .A2(n5438), .A3(n5437), .ZN(n3485) );
  NAND2_X1 U4805 ( .A1(n5466), .A2(b[20]), .ZN(n5363) );
  INV_X1 U4806 ( .A(n5415), .ZN(n5407) );
  INV_X1 U4810 ( .A(n5368), .ZN(n5367) );
  NOR2_X2 U4811 ( .A1(n5336), .A2(n5221), .ZN(n5339) );
  NAND2_X1 U4812 ( .A1(n5525), .A2(b[22]), .ZN(n3271) );
  INV_X1 U4813 ( .A(n5235), .ZN(n3443) );
  INV_X1 U4815 ( .A(n5208), .ZN(n5211) );
  NOR2_X2 U4816 ( .A1(n5348), .A2(n5347), .ZN(n5491) );
  INV_X1 U4817 ( .A(n5488), .ZN(n5485) );
  NAND2_X1 U4818 ( .A1(n5488), .A2(n5484), .ZN(n5486) );
  AOI22_X1 U4819 ( .A1(n5948), .A2(b[23]), .B1(n6043), .B2(b[22]), .ZN(n5949)
         );
  INV_X1 U4820 ( .A(n5894), .ZN(n5896) );
  NAND3_X1 U4821 ( .A1(n6040), .A2(n566), .A3(n6038), .ZN(n6045) );
  OAI21_X1 U4822 ( .B1(n426), .B2(n4096), .A(n4100), .ZN(n4098) );
  INV_X1 U4823 ( .A(n4164), .ZN(n4169) );
  NOR2_X1 U4824 ( .A1(n3984), .A2(n1175), .ZN(n3847) );
  NAND2_X1 U4825 ( .A1(n3984), .A2(n1175), .ZN(n3846) );
  NOR2_X1 U4827 ( .A1(n6376), .A2(n2938), .ZN(n3007) );
  INV_X1 U4828 ( .A(n4978), .ZN(n4980) );
  INV_X1 U4829 ( .A(n5522), .ZN(n5520) );
  OAI21_X1 U4830 ( .B1(n6074), .B2(n6077), .A(n6075), .ZN(n5938) );
  INV_X1 U4831 ( .A(n4142), .ZN(n4140) );
  NAND2_X1 U4832 ( .A1(n4598), .A2(n4219), .ZN(n4110) );
  NAND2_X1 U4834 ( .A1(n5693), .A2(n5688), .ZN(n5690) );
  NOR3_X1 U4835 ( .A1(n3416), .A2(n903), .A3(n6505), .ZN(n3414) );
  INV_X1 U4836 ( .A(n5858), .ZN(n3719) );
  OAI21_X1 U4837 ( .B1(n5600), .B2(n1355), .A(n6661), .ZN(n5605) );
  NAND2_X1 U4838 ( .A1(n1023), .A2(n5332), .ZN(n5333) );
  NAND2_X2 U4839 ( .A1(n6509), .A2(n2711), .ZN(n6009) );
  AOI21_X1 U4841 ( .B1(n6124), .B2(n6123), .A(n6122), .ZN(n6125) );
  AOI21_X1 U4842 ( .B1(n6114), .B2(n6113), .A(n6112), .ZN(n6128) );
  NOR2_X1 U4843 ( .A1(n5827), .A2(n5828), .ZN(n5831) );
  NOR2_X1 U4845 ( .A1(n3387), .A2(n5861), .ZN(n3721) );
  AOI22_X1 U4846 ( .A1(n3718), .A2(n3387), .B1(n3717), .B2(n5858), .ZN(n3716)
         );
  INV_X1 U4847 ( .A(n5861), .ZN(n3717) );
  NAND2_X1 U4848 ( .A1(n3718), .A2(n5850), .ZN(n3715) );
  NOR2_X1 U4853 ( .A1(n6006), .A2(n5998), .ZN(n6008) );
  OAI21_X1 U4854 ( .B1(n6006), .B2(n1314), .A(n6004), .ZN(n6007) );
  AOI21_X1 U4855 ( .B1(n6003), .B2(n6072), .A(n6002), .ZN(n6004) );
  INV_X1 U4857 ( .A(n5878), .ZN(n5879) );
  OAI21_X1 U4858 ( .B1(n5995), .B2(n5583), .A(n5577), .ZN(n5586) );
  NAND2_X1 U4861 ( .A1(n6108), .A2(n6113), .ZN(n6137) );
  XNOR2_X1 U4863 ( .A(n5646), .B(n5645), .ZN(\d[2] ) );
  INV_X1 U4864 ( .A(n5644), .ZN(n5645) );
  XNOR2_X1 U4865 ( .A(n5654), .B(n5653), .ZN(\d[4]_BAR ) );
  AOI21_X1 U4866 ( .B1(n5652), .B2(n6098), .A(n5651), .ZN(n5653) );
  XNOR2_X1 U4867 ( .A(n5660), .B(n5661), .ZN(\d[5]_BAR ) );
  XNOR2_X1 U4868 ( .A(n5658), .B(n5659), .ZN(n5661) );
  XNOR2_X1 U4869 ( .A(n5669), .B(n5668), .ZN(\d[7]_BAR ) );
  AOI21_X1 U4870 ( .B1(n688), .B2(n422), .A(n5666), .ZN(n5668) );
  OAI21_X1 U4871 ( .B1(n5677), .B2(n5674), .A(n5673), .ZN(\d[8]_BAR ) );
  INV_X1 U4872 ( .A(n421), .ZN(n5674) );
  XNOR2_X1 U4873 ( .A(n5680), .B(n5679), .ZN(\d[9]_BAR ) );
  XNOR2_X1 U4874 ( .A(n5702), .B(n5701), .ZN(\d[11]_BAR ) );
  NAND2_X1 U4875 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  XNOR2_X1 U4876 ( .A(n5705), .B(n5706), .ZN(\d[12]_BAR ) );
  OAI21_X1 U4878 ( .B1(n5803), .B2(n5802), .A(n5801), .ZN(\d[20] ) );
  NAND2_X1 U4881 ( .A1(n5811), .A2(n5812), .ZN(n5810) );
  INV_X8 U4882 ( .A(b[3]), .ZN(n3538) );
  XOR2_X2 U4883 ( .A(b[19]), .B(a[9]), .Z(n2702) );
  XOR2_X2 U4885 ( .A(a[11]), .B(b[13]), .Z(n2704) );
  XOR2_X2 U4886 ( .A(a[5]), .B(b[15]), .Z(n2709) );
  XOR2_X2 U4887 ( .A(b[17]), .B(a[9]), .Z(n2710) );
  XOR2_X2 U4888 ( .A(a[7]), .B(b[21]), .Z(n2713) );
  INV_X4 U4889 ( .A(n4522), .ZN(n2774) );
  XOR2_X2 U4890 ( .A(a[19]), .B(b[5]), .Z(n2717) );
  XOR2_X2 U4891 ( .A(a[7]), .B(b[9]), .Z(n2718) );
  XOR2_X2 U4893 ( .A(a[11]), .B(b[3]), .Z(n2723) );
  XNOR2_X2 U4895 ( .A(n5432), .B(n5540), .ZN(n2725) );
  XOR2_X2 U4896 ( .A(a[3]), .B(b[22]), .Z(n2726) );
  XOR2_X2 U4897 ( .A(a[17]), .B(b[9]), .Z(n2727) );
  XOR2_X2 U4898 ( .A(a[17]), .B(b[7]), .Z(n2729) );
  XOR2_X2 U4900 ( .A(a[13]), .B(b[4]), .Z(n2732) );
  INV_X4 U4902 ( .A(n3359), .ZN(n3476) );
  XOR2_X2 U4904 ( .A(a[19]), .B(b[6]), .Z(n2738) );
  XOR2_X2 U4905 ( .A(b[11]), .B(a[19]), .Z(n2739) );
  AND3_X1 U4906 ( .A1(n3639), .A2(a[7]), .A3(b[15]), .ZN(n2740) );
  XOR2_X2 U4907 ( .A(a[15]), .B(b[7]), .Z(n2745) );
  INV_X1 U4908 ( .A(n4599), .ZN(n3607) );
  AND2_X4 U4909 ( .A1(n5919), .A2(n3392), .ZN(n2747) );
  NOR2_X1 U4911 ( .A1(n4873), .A2(n3835), .ZN(n4783) );
  NOR2_X4 U4912 ( .A1(a[22]), .A2(a[21]), .ZN(n4845) );
  NOR2_X2 U4914 ( .A1(n4921), .A2(n4920), .ZN(n5025) );
  OAI21_X2 U4915 ( .B1(n3399), .B2(n3402), .A(n3311), .ZN(n2754) );
  NAND3_X2 U4916 ( .A1(n2759), .A2(n2760), .A3(n5046), .ZN(n5144) );
  NAND2_X2 U4917 ( .A1(n5048), .A2(n5047), .ZN(n2760) );
  NOR2_X2 U4918 ( .A1(n2762), .A2(n5045), .ZN(n2761) );
  INV_X2 U4919 ( .A(n5050), .ZN(n2762) );
  NAND2_X2 U4920 ( .A1(n2764), .A2(n5046), .ZN(n2763) );
  NOR2_X2 U4924 ( .A1(n5394), .A2(n3359), .ZN(n2768) );
  INV_X2 U4925 ( .A(n5926), .ZN(n5394) );
  NAND2_X2 U4926 ( .A1(n483), .A2(n5011), .ZN(n2770) );
  AOI21_X2 U4927 ( .B1(n4957), .B2(n4956), .A(n4955), .ZN(n5011) );
  INV_X2 U4928 ( .A(n4552), .ZN(n2772) );
  OAI21_X1 U4930 ( .B1(n2740), .B2(n4933), .A(n4533), .ZN(n2777) );
  NAND2_X2 U4933 ( .A1(n2781), .A2(n2780), .ZN(n2778) );
  NAND2_X2 U4934 ( .A1(n2779), .A2(n5837), .ZN(n3390) );
  NAND2_X2 U4935 ( .A1(n1099), .A2(n5842), .ZN(n5837) );
  INV_X2 U4936 ( .A(n5624), .ZN(n2782) );
  NAND2_X2 U4937 ( .A1(n3663), .A2(n5375), .ZN(n2822) );
  NAND3_X2 U4938 ( .A1(n3663), .A2(n5375), .A3(n5623), .ZN(n2784) );
  INV_X2 U4939 ( .A(n5623), .ZN(n2786) );
  NOR2_X4 U4940 ( .A1(n3321), .A2(n4971), .ZN(n5842) );
  NOR2_X2 U4942 ( .A1(n3177), .A2(n3175), .ZN(n2793) );
  OAI22_X2 U4943 ( .A1(n5074), .A2(b[12]), .B1(n440), .B2(n5277), .ZN(n2794)
         );
  NAND2_X2 U4944 ( .A1(n1326), .A2(n2704), .ZN(n2795) );
  NOR2_X2 U4946 ( .A1(n2799), .A2(n5088), .ZN(n2798) );
  NOR2_X1 U4947 ( .A1(n4703), .A2(n3598), .ZN(n2800) );
  AOI22_X2 U4949 ( .A1(n5900), .A2(b[8]), .B1(n3342), .B2(n435), .ZN(n4947) );
  NAND2_X2 U4951 ( .A1(n3216), .A2(n4496), .ZN(n4555) );
  NAND2_X2 U4952 ( .A1(n2807), .A2(n5601), .ZN(n5608) );
  NOR2_X2 U4953 ( .A1(n5993), .A2(n5992), .ZN(\d[37]_BAR ) );
  NAND2_X2 U4954 ( .A1(n2809), .A2(n3943), .ZN(n4055) );
  NOR2_X2 U4955 ( .A1(n2809), .A2(n3943), .ZN(n4060) );
  NAND2_X2 U4956 ( .A1(n5353), .A2(n2810), .ZN(n2846) );
  NAND2_X2 U4957 ( .A1(n2815), .A2(n2816), .ZN(n2811) );
  NAND2_X2 U4959 ( .A1(n6043), .A2(b[14]), .ZN(n2815) );
  NAND2_X2 U4960 ( .A1(n3142), .A2(n5293), .ZN(n2816) );
  NAND2_X2 U4961 ( .A1(n5476), .A2(n984), .ZN(n2817) );
  NAND2_X1 U4962 ( .A1(n3351), .A2(n5105), .ZN(n3272) );
  NOR2_X2 U4964 ( .A1(n2822), .A2(n3725), .ZN(n6013) );
  NAND2_X2 U4965 ( .A1(n4950), .A2(n4951), .ZN(n5023) );
  INV_X4 U4967 ( .A(n4933), .ZN(n2828) );
  INV_X8 U4968 ( .A(n2829), .ZN(n2830) );
  NAND2_X2 U4970 ( .A1(n2831), .A2(n3288), .ZN(n5772) );
  NOR3_X2 U4971 ( .A1(n2832), .A2(n3391), .A3(n4971), .ZN(n5850) );
  INV_X2 U4972 ( .A(n5919), .ZN(n3391) );
  NAND2_X2 U4973 ( .A1(n5887), .A2(n289), .ZN(n4971) );
  AOI21_X1 U4974 ( .B1(n3098), .B2(n3353), .A(n3428), .ZN(n2832) );
  INV_X2 U4975 ( .A(n4719), .ZN(n4721) );
  INV_X8 U4977 ( .A(n2828), .ZN(n3405) );
  NAND2_X2 U4980 ( .A1(n3605), .A2(n3606), .ZN(n2841) );
  INV_X2 U4982 ( .A(n4603), .ZN(n2842) );
  NOR2_X2 U4983 ( .A1(n3573), .A2(n4602), .ZN(n4603) );
  NAND2_X2 U4984 ( .A1(n2843), .A2(n2845), .ZN(n2844) );
  NOR2_X1 U4987 ( .A1(b[17]), .A2(n4940), .ZN(n2850) );
  AOI21_X2 U4988 ( .B1(n6111), .B2(n2908), .A(n882), .ZN(n2851) );
  NAND3_X2 U4990 ( .A1(n1042), .A2(n5173), .A3(n5174), .ZN(n2856) );
  NAND2_X2 U4991 ( .A1(n5141), .A2(n5140), .ZN(n5175) );
  BUF_X4 U4992 ( .A(n2932), .Z(n2858) );
  NAND2_X2 U4993 ( .A1(n2860), .A2(n2859), .ZN(n5135) );
  NAND2_X1 U4994 ( .A1(n2932), .A2(n3372), .ZN(n2859) );
  NAND2_X2 U4996 ( .A1(n2867), .A2(n2866), .ZN(n3977) );
  INV_X2 U4997 ( .A(n4634), .ZN(n5757) );
  NAND2_X2 U5000 ( .A1(n2858), .A2(n2875), .ZN(n2873) );
  AOI21_X2 U5001 ( .B1(n5340), .B2(n2858), .A(n2875), .ZN(n2874) );
  INV_X2 U5002 ( .A(n5450), .ZN(n2875) );
  NAND2_X2 U5005 ( .A1(n6072), .A2(n6071), .ZN(n6086) );
  NOR2_X2 U5006 ( .A1(n5612), .A2(n369), .ZN(n6072) );
  AOI21_X2 U5007 ( .B1(n6526), .B2(n259), .A(n5394), .ZN(n6071) );
  NOR2_X4 U5012 ( .A1(n2830), .A2(n4988), .ZN(n3532) );
  NAND2_X2 U5013 ( .A1(n5098), .A2(n5097), .ZN(n2879) );
  AOI22_X1 U5014 ( .A1(n4780), .A2(n3313), .B1(n4779), .B2(n1440), .ZN(n2880)
         );
  INV_X1 U5016 ( .A(n4686), .ZN(n2886) );
  NOR2_X1 U5017 ( .A1(n1018), .A2(n4643), .ZN(n4647) );
  INV_X1 U5019 ( .A(n5628), .ZN(n5969) );
  NOR2_X2 U5021 ( .A1(n3105), .A2(n5603), .ZN(n5604) );
  NAND2_X1 U5022 ( .A1(n3567), .A2(n5621), .ZN(n5624) );
  NOR2_X4 U5024 ( .A1(n3111), .A2(n5233), .ZN(n5234) );
  AOI21_X1 U5025 ( .B1(n3870), .B2(n6328), .A(n5952), .ZN(n4815) );
  NAND2_X2 U5026 ( .A1(n6095), .A2(n2892), .ZN(n2893) );
  NAND2_X2 U5027 ( .A1(n2893), .A2(n2894), .ZN(\d[25] ) );
  INV_X1 U5029 ( .A(n6095), .ZN(n6094) );
  NAND2_X1 U5030 ( .A1(n5161), .A2(n5162), .ZN(n5163) );
  INV_X1 U5031 ( .A(n5723), .ZN(n5724) );
  OAI21_X1 U5032 ( .B1(n438), .B2(n5717), .A(n2294), .ZN(n5719) );
  NOR2_X1 U5034 ( .A1(n4002), .A2(n3798), .ZN(n3797) );
  NAND2_X2 U5036 ( .A1(n6199), .A2(n3155), .ZN(n2900) );
  NOR2_X1 U5038 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  NOR2_X1 U5039 ( .A1(n5583), .A2(n6000), .ZN(n5584) );
  NAND3_X1 U5040 ( .A1(n5582), .A2(n6000), .A3(n5995), .ZN(n5591) );
  INV_X1 U5041 ( .A(n6000), .ZN(n5871) );
  INV_X1 U5042 ( .A(n5602), .ZN(n5603) );
  NAND2_X1 U5045 ( .A1(n5767), .A2(n5727), .ZN(n5746) );
  NOR2_X1 U5046 ( .A1(n5634), .A2(n1355), .ZN(n5631) );
  INV_X1 U5047 ( .A(n4639), .ZN(n4641) );
  INV_X1 U5049 ( .A(n5377), .ZN(n5378) );
  AOI22_X1 U5050 ( .A1(n3007), .A2(n2937), .B1(n6447), .B2(n6376), .ZN(n3001)
         );
  NOR2_X4 U5055 ( .A1(n5362), .A2(n5361), .ZN(n5459) );
  AOI22_X2 U5057 ( .A1(n3308), .A2(n4349), .B1(n4351), .B2(n4350), .ZN(n2906)
         );
  NAND2_X4 U5058 ( .A1(a[17]), .A2(a[18]), .ZN(n2911) );
  INV_X8 U5060 ( .A(a[18]), .ZN(n2910) );
  NAND2_X1 U5061 ( .A1(n5360), .A2(a[23]), .ZN(n5530) );
  NAND2_X1 U5062 ( .A1(n5235), .A2(n5360), .ZN(n3310) );
  NOR2_X1 U5063 ( .A1(n5360), .A2(n4601), .ZN(n3432) );
  NAND2_X1 U5064 ( .A1(n6185), .A2(n2603), .ZN(n4129) );
  NOR2_X1 U5065 ( .A1(n2603), .A2(n6616), .ZN(n3992) );
  NOR3_X2 U5067 ( .A1(n5396), .A2(n2915), .A3(n2914), .ZN(n5420) );
  NAND2_X2 U5070 ( .A1(n3424), .A2(n3464), .ZN(n3423) );
  XNOR2_X2 U5072 ( .A(n4793), .B(n4953), .ZN(n4961) );
  NAND2_X2 U5080 ( .A1(n4012), .A2(n4013), .ZN(n2927) );
  BUF_X4 U5081 ( .A(n2929), .Z(n2928) );
  NAND2_X2 U5082 ( .A1(n3004), .A2(n3001), .ZN(n4631) );
  AOI21_X2 U5083 ( .B1(n1043), .B2(n3570), .A(n4521), .ZN(n4575) );
  NOR2_X2 U5084 ( .A1(n4572), .A2(n4574), .ZN(n2930) );
  INV_X4 U5085 ( .A(n2933), .ZN(n5381) );
  NAND2_X2 U5086 ( .A1(n5382), .A2(n5625), .ZN(n2936) );
  NOR2_X2 U5087 ( .A1(n2935), .A2(n2934), .ZN(n5385) );
  NAND2_X2 U5088 ( .A1(n5625), .A2(n2747), .ZN(n2934) );
  INV_X2 U5089 ( .A(n5382), .ZN(n2935) );
  AOI22_X1 U5090 ( .A1(n2936), .A2(n5390), .B1(n5620), .B2(n3392), .ZN(n5391)
         );
  INV_X4 U5091 ( .A(n2939), .ZN(n2938) );
  NAND2_X2 U5092 ( .A1(n2941), .A2(n2940), .ZN(n4553) );
  NAND3_X2 U5093 ( .A1(n2944), .A2(n2943), .A3(n2942), .ZN(n2941) );
  INV_X2 U5094 ( .A(n2946), .ZN(n2944) );
  NAND2_X2 U5097 ( .A1(n3170), .A2(n6325), .ZN(n2948) );
  AOI21_X2 U5098 ( .B1(n3289), .B2(n3288), .A(n3287), .ZN(n2951) );
  NOR2_X2 U5099 ( .A1(n1909), .A2(n4315), .ZN(n2952) );
  NAND2_X1 U5101 ( .A1(a[19]), .A2(n2954), .ZN(n5522) );
  NAND2_X2 U5103 ( .A1(n2963), .A2(n2959), .ZN(n3541) );
  INV_X2 U5107 ( .A(n4759), .ZN(n2964) );
  BUF_X4 U5108 ( .A(n5793), .Z(n2970) );
  NAND2_X2 U5109 ( .A1(n1046), .A2(n3914), .ZN(n2975) );
  BUF_X4 U5110 ( .A(n343), .Z(n2976) );
  NOR2_X2 U5112 ( .A1(n6008), .A2(n6007), .ZN(n2981) );
  INV_X2 U5113 ( .A(n3612), .ZN(n2982) );
  BUF_X4 U5115 ( .A(n5665), .Z(n2984) );
  AOI21_X2 U5116 ( .B1(n4428), .B2(n3562), .A(n4427), .ZN(n4442) );
  BUF_X4 U5117 ( .A(n1059), .Z(n2985) );
  OAI21_X2 U5118 ( .B1(n4984), .B2(n4983), .A(n997), .ZN(n4985) );
  AOI21_X2 U5120 ( .B1(n4379), .B2(n4378), .A(n2991), .ZN(n2990) );
  NOR2_X2 U5123 ( .A1(n2992), .A2(n4018), .ZN(n4379) );
  AOI22_X2 U5124 ( .A1(n397), .A2(n4016), .B1(n4017), .B2(n2994), .ZN(n3495)
         );
  NAND2_X2 U5125 ( .A1(n4954), .A2(n4956), .ZN(n4793) );
  NAND2_X2 U5126 ( .A1(n4786), .A2(n3000), .ZN(n4956) );
  NAND2_X2 U5127 ( .A1(n2999), .A2(n4785), .ZN(n4954) );
  INV_X2 U5128 ( .A(n3000), .ZN(n2999) );
  AOI21_X2 U5129 ( .B1(n4782), .B2(n3203), .A(n4783), .ZN(n3000) );
  NAND2_X2 U5132 ( .A1(n3006), .A2(n3005), .ZN(n3004) );
  INV_X2 U5133 ( .A(n3007), .ZN(n3006) );
  INV_X2 U5134 ( .A(n4008), .ZN(n3009) );
  AOI22_X2 U5136 ( .A1(n3870), .A2(n3011), .B1(n5041), .B2(b[5]), .ZN(n3923)
         );
  NAND2_X2 U5138 ( .A1(n3371), .A2(n5315), .ZN(n3012) );
  AOI22_X2 U5139 ( .A1(n4654), .A2(n3014), .B1(n800), .B2(n3013), .ZN(n4736)
         );
  AOI22_X2 U5142 ( .A1(n4625), .A2(n6570), .B1(n1040), .B2(n4623), .ZN(n4654)
         );
  AOI21_X2 U5143 ( .B1(n975), .B2(n3020), .A(n3018), .ZN(n4384) );
  NAND2_X2 U5144 ( .A1(n3019), .A2(n6528), .ZN(n3018) );
  NAND2_X2 U5145 ( .A1(n4337), .A2(b[16]), .ZN(n3019) );
  INV_X8 U5146 ( .A(a[19]), .ZN(n4026) );
  NAND2_X2 U5147 ( .A1(n3472), .A2(n3242), .ZN(n3028) );
  NAND2_X2 U5149 ( .A1(n3031), .A2(n3831), .ZN(n3030) );
  XNOR2_X1 U5150 ( .A(n678), .B(n4259), .ZN(n4265) );
  NAND2_X2 U5151 ( .A1(n3320), .A2(n4211), .ZN(n3036) );
  INV_X2 U5152 ( .A(n4250), .ZN(n3037) );
  NAND2_X2 U5153 ( .A1(n3040), .A2(n3039), .ZN(n3038) );
  NAND3_X2 U5154 ( .A1(n4211), .A2(n4249), .A3(n3320), .ZN(n3039) );
  OAI21_X2 U5155 ( .B1(n4466), .B2(n3349), .A(n579), .ZN(n3041) );
  INV_X4 U5156 ( .A(n3043), .ZN(n4042) );
  NAND2_X1 U5158 ( .A1(n3045), .A2(n4933), .ZN(n3044) );
  INV_X2 U5159 ( .A(n3960), .ZN(n3045) );
  NAND2_X2 U5160 ( .A1(n3047), .A2(n3617), .ZN(n3046) );
  INV_X2 U5161 ( .A(n3961), .ZN(n3047) );
  INV_X2 U5162 ( .A(n3962), .ZN(n3048) );
  NOR2_X2 U5164 ( .A1(n4999), .A2(b[11]), .ZN(n3055) );
  INV_X2 U5167 ( .A(n4471), .ZN(n3060) );
  NAND2_X2 U5171 ( .A1(n3556), .A2(n4824), .ZN(n3066) );
  INV_X2 U5174 ( .A(n4344), .ZN(n4343) );
  NAND2_X2 U5175 ( .A1(n3072), .A2(n3071), .ZN(n4344) );
  XNOR2_X2 U5176 ( .A(b[18]), .B(a[7]), .ZN(n3080) );
  NAND2_X2 U5177 ( .A1(n4705), .A2(b[13]), .ZN(n3081) );
  NAND2_X2 U5178 ( .A1(n2726), .A2(n1059), .ZN(n3084) );
  NAND2_X2 U5179 ( .A1(n4467), .A2(n4468), .ZN(n3087) );
  NAND2_X2 U5180 ( .A1(n4458), .A2(n4459), .ZN(n4468) );
  NAND3_X2 U5181 ( .A1(n5011), .A2(n484), .A3(n808), .ZN(n3091) );
  NAND2_X2 U5182 ( .A1(n3669), .A2(n4958), .ZN(n3092) );
  NAND2_X1 U5183 ( .A1(n5092), .A2(n437), .ZN(n3578) );
  NOR2_X1 U5184 ( .A1(n5092), .A2(n437), .ZN(n3579) );
  BUF_X4 U5186 ( .A(n4637), .Z(n3097) );
  INV_X2 U5187 ( .A(n5850), .ZN(n3102) );
  OAI21_X1 U5188 ( .B1(n5850), .B2(n3387), .A(n3099), .ZN(n3101) );
  NAND3_X2 U5189 ( .A1(n3102), .A2(n3406), .A3(n5856), .ZN(n3100) );
  NAND3_X2 U5190 ( .A1(n3100), .A2(n3101), .A3(n5857), .ZN(\d[30] ) );
  NAND2_X1 U5192 ( .A1(n690), .A2(n432), .ZN(n4966) );
  BUF_X4 U5194 ( .A(n2830), .Z(n3111) );
  NAND2_X2 U5196 ( .A1(n2827), .A2(n4879), .ZN(n3560) );
  INV_X2 U5198 ( .A(n6006), .ZN(n3117) );
  NAND2_X2 U5199 ( .A1(n3120), .A2(n3190), .ZN(n3119) );
  NAND2_X4 U5203 ( .A1(n5860), .A2(n5859), .ZN(n5094) );
  INV_X8 U5204 ( .A(n4933), .ZN(n3617) );
  AOI22_X2 U5206 ( .A1(n3377), .A2(n3378), .B1(n482), .B2(n3379), .ZN(n5037)
         );
  NAND2_X2 U5208 ( .A1(n4372), .A2(n4373), .ZN(n3569) );
  INV_X2 U5209 ( .A(b[17]), .ZN(n3131) );
  BUF_X4 U5210 ( .A(n3317), .Z(n3133) );
  BUF_X4 U5212 ( .A(n5764), .Z(n3135) );
  NOR2_X2 U5215 ( .A1(n3138), .A2(n4985), .ZN(\d[31] ) );
  NAND2_X2 U5217 ( .A1(n3139), .A2(n5810), .ZN(\d[27]_BAR ) );
  NAND2_X2 U5218 ( .A1(n3141), .A2(n3140), .ZN(n3139) );
  INV_X2 U5219 ( .A(n5811), .ZN(n3141) );
  INV_X8 U5220 ( .A(b[21]), .ZN(n5951) );
  BUF_X4 U5221 ( .A(n5477), .Z(n3142) );
  NAND2_X2 U5222 ( .A1(n6131), .A2(n6130), .ZN(n3143) );
  NAND2_X2 U5223 ( .A1(b[13]), .A2(n5900), .ZN(n3144) );
  NAND2_X2 U5224 ( .A1(n5947), .A2(n184), .ZN(n3145) );
  INV_X4 U5226 ( .A(n4885), .ZN(n3252) );
  NOR2_X2 U5227 ( .A1(n3704), .A2(n4595), .ZN(n4596) );
  NAND2_X2 U5228 ( .A1(n6213), .A2(n4332), .ZN(n3146) );
  NAND2_X4 U5229 ( .A1(n3308), .A2(b[0]), .ZN(n4035) );
  NAND2_X2 U5231 ( .A1(n4705), .A2(b[9]), .ZN(n3148) );
  INV_X2 U5233 ( .A(n5700), .ZN(n3151) );
  NAND2_X2 U5234 ( .A1(n3364), .A2(n3363), .ZN(n5700) );
  NOR2_X4 U5235 ( .A1(n506), .A2(a[5]), .ZN(n4504) );
  INV_X4 U5236 ( .A(n3360), .ZN(n5926) );
  NAND2_X4 U5237 ( .A1(n3153), .A2(n3452), .ZN(n5682) );
  BUF_X4 U5238 ( .A(n6134), .Z(n3157) );
  NAND2_X2 U5239 ( .A1(n5356), .A2(n5355), .ZN(n3158) );
  INV_X8 U5240 ( .A(a[0]), .ZN(n4490) );
  OAI211_X1 U5241 ( .C1(n6138), .C2(n6137), .A(n3159), .B(n6136), .ZN(\d[47] )
         );
  BUF_X4 U5242 ( .A(n4940), .Z(n3161) );
  INV_X2 U5243 ( .A(n3790), .ZN(n3418) );
  NAND2_X2 U5244 ( .A1(n3163), .A2(n3162), .ZN(n3790) );
  NAND2_X2 U5245 ( .A1(n5110), .A2(b[0]), .ZN(n3162) );
  BUF_X4 U5246 ( .A(n5999), .Z(n3164) );
  NAND3_X2 U5247 ( .A1(n3390), .A2(n3678), .A3(n5627), .ZN(n3676) );
  BUF_X4 U5249 ( .A(n5707), .Z(n3167) );
  INV_X8 U5250 ( .A(n4010), .ZN(n4408) );
  NOR2_X4 U5252 ( .A1(n4973), .A2(n4974), .ZN(n5808) );
  INV_X2 U5254 ( .A(n3983), .ZN(n3276) );
  NAND2_X2 U5257 ( .A1(n3180), .A2(n3885), .ZN(n3179) );
  NAND2_X2 U5258 ( .A1(n3482), .A2(n3914), .ZN(n3180) );
  INV_X2 U5259 ( .A(n4685), .ZN(n3181) );
  NOR2_X2 U5260 ( .A1(n4597), .A2(n4596), .ZN(n4685) );
  NAND3_X2 U5262 ( .A1(n1046), .A2(n3482), .A3(n3914), .ZN(n3182) );
  NOR2_X2 U5263 ( .A1(n3912), .A2(n3868), .ZN(n3183) );
  NOR2_X2 U5265 ( .A1(n5565), .A2(n1100), .ZN(n3193) );
  NAND2_X2 U5266 ( .A1(n5565), .A2(n1100), .ZN(n3194) );
  NOR2_X2 U5267 ( .A1(n5506), .A2(n5507), .ZN(n5551) );
  AOI22_X2 U5268 ( .A1(n3195), .A2(n416), .B1(n5458), .B2(n5459), .ZN(n5507)
         );
  NAND2_X2 U5270 ( .A1(n6528), .A2(n3431), .ZN(n3556) );
  MUX2_X2 U5273 ( .A(n3431), .B(n4504), .S(b[14]), .Z(n3941) );
  MUX2_X2 U5274 ( .A(n3431), .B(n4504), .S(b[6]), .Z(n4226) );
  NAND2_X2 U5277 ( .A1(n501), .A2(n3369), .ZN(n3368) );
  NAND2_X2 U5278 ( .A1(n4551), .A2(n3510), .ZN(n3215) );
  INV_X1 U5280 ( .A(n3581), .ZN(n4772) );
  NAND2_X2 U5281 ( .A1(n3334), .A2(n5193), .ZN(n5194) );
  NAND2_X2 U5282 ( .A1(n3334), .A2(n5137), .ZN(n5138) );
  NOR2_X2 U5285 ( .A1(n4659), .A2(n945), .ZN(n3223) );
  INV_X2 U5286 ( .A(n3224), .ZN(n4406) );
  OAI21_X2 U5289 ( .B1(n3964), .B2(n3963), .A(n3226), .ZN(n4039) );
  NAND2_X1 U5290 ( .A1(n2744), .A2(n1059), .ZN(n3226) );
  BUF_X4 U5291 ( .A(n5473), .Z(n3230) );
  NAND3_X2 U5292 ( .A1(n3233), .A2(n5843), .A3(n5840), .ZN(n5848) );
  NAND2_X2 U5293 ( .A1(n5838), .A2(n1099), .ZN(n3233) );
  NAND3_X2 U5297 ( .A1(n2736), .A2(n3247), .A3(n3246), .ZN(n3245) );
  INV_X2 U5299 ( .A(n3250), .ZN(n4870) );
  INV_X1 U5300 ( .A(n4539), .ZN(n3253) );
  INV_X2 U5301 ( .A(n4589), .ZN(n3254) );
  INV_X4 U5302 ( .A(n5041), .ZN(n5106) );
  NOR2_X4 U5303 ( .A1(a[13]), .A2(a[11]), .ZN(n3258) );
  NOR2_X4 U5304 ( .A1(a[12]), .A2(a[13]), .ZN(n3259) );
  INV_X2 U5307 ( .A(b[17]), .ZN(n3263) );
  NOR2_X2 U5308 ( .A1(n4858), .A2(n4857), .ZN(n4884) );
  NOR2_X1 U5310 ( .A1(n3269), .A2(n5030), .ZN(n3749) );
  NAND3_X2 U5311 ( .A1(n3280), .A2(n3279), .A3(n3278), .ZN(n3277) );
  NAND3_X2 U5312 ( .A1(n4751), .A2(n4846), .A3(b[5]), .ZN(n3279) );
  INV_X2 U5315 ( .A(n4627), .ZN(n3285) );
  NOR2_X2 U5317 ( .A1(n4292), .A2(n4005), .ZN(n3287) );
  NAND2_X2 U5318 ( .A1(n4292), .A2(n4005), .ZN(n3288) );
  INV_X2 U5319 ( .A(n3642), .ZN(n3293) );
  NAND2_X4 U5323 ( .A1(a[8]), .A2(a[7]), .ZN(n3305) );
  NOR2_X4 U5324 ( .A1(n3305), .A2(a[9]), .ZN(n4794) );
  NAND2_X2 U5325 ( .A1(n3307), .A2(n3306), .ZN(n3695) );
  INV_X4 U5326 ( .A(n3562), .ZN(n3699) );
  INV_X2 U5328 ( .A(n4925), .ZN(n3311) );
  OAI21_X2 U5329 ( .B1(n3416), .B2(n903), .A(n5700), .ZN(n3317) );
  INV_X1 U5330 ( .A(n5808), .ZN(n5841) );
  OAI21_X1 U5333 ( .B1(n3340), .B2(n4630), .A(n4629), .ZN(n3339) );
  NOR2_X2 U5334 ( .A1(n6156), .A2(n3343), .ZN(n4019) );
  MUX2_X2 U5336 ( .A(n5525), .B(n3351), .S(n1896), .Z(n5528) );
  NOR2_X1 U5338 ( .A1(n5853), .A2(n3354), .ZN(n5856) );
  INV_X2 U5341 ( .A(n4288), .ZN(n3357) );
  OAI22_X2 U5342 ( .A1(n5847), .A2(n5846), .B1(n5848), .B2(n5849), .ZN(\d[28] ) );
  NAND2_X2 U5343 ( .A1(n3362), .A2(n2294), .ZN(n3361) );
  INV_X2 U5344 ( .A(n4266), .ZN(n3363) );
  NAND2_X2 U5345 ( .A1(n5681), .A2(n5685), .ZN(n3365) );
  NOR2_X4 U5346 ( .A1(n5682), .A2(n3366), .ZN(n3416) );
  NOR2_X2 U5347 ( .A1(n5681), .A2(n5685), .ZN(n3366) );
  OAI21_X2 U5348 ( .B1(n3985), .B2(n3847), .A(n3846), .ZN(n4315) );
  NAND3_X1 U5349 ( .A1(n4415), .A2(n3369), .A3(n3870), .ZN(n4358) );
  NAND2_X2 U5350 ( .A1(n3374), .A2(n3373), .ZN(n4781) );
  NAND2_X2 U5351 ( .A1(n2858), .A2(n3020), .ZN(n3373) );
  NAND2_X2 U5352 ( .A1(n984), .A2(n512), .ZN(n3381) );
  NAND2_X2 U5353 ( .A1(n5951), .A2(n3326), .ZN(n3601) );
  NAND2_X2 U5355 ( .A1(n3407), .A2(n3551), .ZN(n3387) );
  NOR2_X2 U5356 ( .A1(n3388), .A2(n5850), .ZN(n4984) );
  NOR2_X2 U5357 ( .A1(n5624), .A2(n3726), .ZN(n5623) );
  INV_X4 U5358 ( .A(n4887), .ZN(n4590) );
  NAND3_X1 U5360 ( .A1(n3394), .A2(a[13]), .A3(b[5]), .ZN(n4357) );
  NOR2_X4 U5361 ( .A1(n908), .A2(n5733), .ZN(n5729) );
  NAND2_X2 U5362 ( .A1(n3401), .A2(n3400), .ZN(n3399) );
  NAND2_X2 U5363 ( .A1(n3020), .A2(n5076), .ZN(n3400) );
  INV_X2 U5365 ( .A(n3789), .ZN(n3417) );
  AOI21_X2 U5366 ( .B1(n3420), .B2(n3422), .A(n3419), .ZN(n3842) );
  NOR3_X2 U5367 ( .A1(n3789), .A2(n3422), .A3(n3790), .ZN(n3419) );
  INV_X2 U5368 ( .A(n3824), .ZN(n3422) );
  NAND2_X2 U5369 ( .A1(n4272), .A2(n3425), .ZN(n3424) );
  INV_X2 U5370 ( .A(n4271), .ZN(n3425) );
  NOR2_X2 U5371 ( .A1(n3699), .A2(n4943), .ZN(n5015) );
  INV_X4 U5373 ( .A(n5918), .ZN(n5887) );
  INV_X2 U5374 ( .A(n4550), .ZN(n3429) );
  NOR2_X2 U5375 ( .A1(n3614), .A2(b[18]), .ZN(n3433) );
  NOR2_X2 U5379 ( .A1(n3443), .A2(n5410), .ZN(n5517) );
  NAND3_X1 U5380 ( .A1(n3020), .A2(a[19]), .A3(n3562), .ZN(n5146) );
  INV_X2 U5381 ( .A(n3444), .ZN(n5468) );
  MUX2_X2 U5382 ( .A(n3445), .B(n5235), .S(n5951), .Z(n3444) );
  INV_X2 U5383 ( .A(n5466), .ZN(n3445) );
  INV_X2 U5384 ( .A(n3622), .ZN(n3451) );
  NOR2_X4 U5385 ( .A1(n3722), .A2(n5672), .ZN(n5678) );
  NAND2_X2 U5386 ( .A1(n3455), .A2(n185), .ZN(n3454) );
  NOR2_X2 U5387 ( .A1(n4187), .A2(n4182), .ZN(n3455) );
  NAND3_X2 U5390 ( .A1(n4230), .A2(n4229), .A3(n4187), .ZN(n3459) );
  BUF_X4 U5391 ( .A(n5794), .Z(n3460) );
  INV_X4 U5392 ( .A(n4312), .ZN(n3461) );
  INV_X2 U5393 ( .A(n3466), .ZN(n5858) );
  OAI21_X2 U5394 ( .B1(n3497), .B2(n5206), .A(n5215), .ZN(n3471) );
  INV_X2 U5395 ( .A(n3921), .ZN(n3475) );
  NOR2_X2 U5398 ( .A1(n3575), .A2(n4919), .ZN(n4891) );
  INV_X2 U5400 ( .A(n5448), .ZN(n5462) );
  INV_X2 U5401 ( .A(n3487), .ZN(n3486) );
  NAND2_X2 U5403 ( .A1(n3490), .A2(n3489), .ZN(n5425) );
  NAND2_X1 U5404 ( .A1(n760), .A2(b[23]), .ZN(n3489) );
  AOI21_X2 U5409 ( .B1(n4454), .B2(n3495), .A(n3737), .ZN(n4459) );
  NOR2_X1 U5410 ( .A1(n3369), .A2(b[6]), .ZN(n4013) );
  INV_X2 U5411 ( .A(n5216), .ZN(n3497) );
  NAND3_X2 U5412 ( .A1(n3499), .A2(n5217), .A3(n5216), .ZN(n3498) );
  XOR2_X2 U5415 ( .A(a[16]), .B(a[15]), .Z(n3506) );
  INV_X2 U5416 ( .A(n4377), .ZN(n3508) );
  INV_X1 U5417 ( .A(n4528), .ZN(n4640) );
  XNOR2_X1 U5418 ( .A(n5663), .B(n688), .ZN(\d[6]_BAR ) );
  INV_X8 U5421 ( .A(n3513), .ZN(n6035) );
  NAND2_X2 U5422 ( .A1(n3515), .A2(n3514), .ZN(n5232) );
  INV_X4 U5423 ( .A(n3518), .ZN(n5290) );
  NAND2_X2 U5424 ( .A1(n3518), .A2(n5289), .ZN(n3558) );
  NAND2_X2 U5426 ( .A1(n4120), .A2(n6528), .ZN(n4141) );
  INV_X8 U5427 ( .A(n4752), .ZN(n5900) );
  BUF_X4 U5429 ( .A(n3520), .Z(n3519) );
  OAI21_X1 U5430 ( .B1(n5829), .B2(n5828), .A(n3519), .ZN(n5830) );
  NAND2_X2 U5431 ( .A1(n3530), .A2(n5048), .ZN(n3528) );
  INV_X2 U5433 ( .A(n3534), .ZN(n5710) );
  NOR2_X2 U5434 ( .A1(n6589), .A2(n4355), .ZN(n4356) );
  XNOR2_X2 U5436 ( .A(n3541), .B(n4707), .ZN(n4738) );
  NOR2_X2 U5437 ( .A1(n3544), .A2(n3543), .ZN(n3542) );
  NOR2_X2 U5439 ( .A1(n2725), .A2(n5574), .ZN(n5914) );
  NAND2_X2 U5440 ( .A1(n3766), .A2(n5415), .ZN(n5417) );
  NAND2_X2 U5441 ( .A1(n3549), .A2(n5422), .ZN(n5415) );
  INV_X2 U5442 ( .A(n1015), .ZN(n3552) );
  INV_X2 U5443 ( .A(n5375), .ZN(n5845) );
  AOI21_X2 U5444 ( .B1(n326), .B2(n4235), .A(n3998), .ZN(n4284) );
  NAND3_X2 U5445 ( .A1(n3998), .A2(n326), .A3(n4235), .ZN(n3582) );
  NAND2_X2 U5447 ( .A1(n2628), .A2(n2627), .ZN(n3559) );
  INV_X8 U5448 ( .A(b[13]), .ZN(n4614) );
  NAND2_X2 U5449 ( .A1(n3566), .A2(n3565), .ZN(n4383) );
  NAND2_X2 U5450 ( .A1(b[15]), .A2(n4506), .ZN(n3565) );
  OAI21_X2 U5451 ( .B1(n4029), .B2(n4028), .A(n3618), .ZN(n4032) );
  INV_X4 U5452 ( .A(n3567), .ZN(n5620) );
  INV_X2 U5454 ( .A(n3582), .ZN(n4283) );
  BUF_X4 U5455 ( .A(n908), .Z(n3590) );
  NAND2_X2 U5457 ( .A1(n3601), .A2(n3600), .ZN(n4930) );
  NAND2_X2 U5458 ( .A1(n4089), .A2(n6528), .ZN(n4166) );
  AOI21_X2 U5459 ( .B1(n4226), .B2(n6558), .A(n4225), .ZN(n4257) );
  AOI22_X2 U5460 ( .A1(n4492), .A2(b[17]), .B1(n6515), .B2(a[3]), .ZN(n3610)
         );
  MUX2_X2 U5461 ( .A(n4600), .B(n4601), .S(b[2]), .Z(n4165) );
  MUX2_X2 U5463 ( .A(n3614), .B(n4601), .S(b[8]), .Z(n3799) );
  NAND2_X2 U5465 ( .A1(n3562), .A2(n2733), .ZN(n3618) );
  INV_X2 U5467 ( .A(n5044), .ZN(n3632) );
  NAND2_X2 U5468 ( .A1(n3637), .A2(n3635), .ZN(n3633) );
  INV_X2 U5469 ( .A(a[9]), .ZN(n3639) );
  NOR2_X2 U5470 ( .A1(a[9]), .A2(b[23]), .ZN(n3636) );
  INV_X2 U5471 ( .A(a[9]), .ZN(n3638) );
  NAND2_X2 U5474 ( .A1(n3884), .A2(n3883), .ZN(n3914) );
  NAND2_X2 U5475 ( .A1(n3651), .A2(n3649), .ZN(n3885) );
  XNOR2_X2 U5476 ( .A(n4195), .B(n6337), .ZN(n3656) );
  NAND2_X2 U5478 ( .A1(n5351), .A2(n5349), .ZN(n3660) );
  INV_X2 U5479 ( .A(n4293), .ZN(n4292) );
  NAND3_X2 U5484 ( .A1(n344), .A2(n5922), .A3(n6350), .ZN(n5313) );
  NAND2_X4 U5486 ( .A1(a[2]), .A2(a[1]), .ZN(n3671) );
  INV_X2 U5487 ( .A(n4891), .ZN(n5026) );
  NAND2_X2 U5489 ( .A1(n3677), .A2(n3676), .ZN(\d[34] ) );
  BUF_X4 U5490 ( .A(n5860), .Z(n3679) );
  AOI22_X2 U5491 ( .A1(n4208), .A2(n4209), .B1(n397), .B2(n4207), .ZN(n4250)
         );
  NAND2_X2 U5492 ( .A1(n3681), .A2(n5990), .ZN(n5992) );
  INV_X2 U5493 ( .A(n5991), .ZN(n3682) );
  INV_X8 U5496 ( .A(a[7]), .ZN(n4689) );
  NAND3_X2 U5497 ( .A1(n5593), .A2(n5595), .A3(n5594), .ZN(\d[43] ) );
  INV_X8 U5498 ( .A(a[9]), .ZN(n3684) );
  INV_X2 U5500 ( .A(n4878), .ZN(n3687) );
  NOR2_X1 U5501 ( .A1(n2705), .A2(n5928), .ZN(n3771) );
  NAND2_X4 U5503 ( .A1(n5070), .A2(a[19]), .ZN(n5180) );
  NOR2_X4 U5504 ( .A1(a[18]), .A2(a[17]), .ZN(n5070) );
  INV_X2 U5506 ( .A(n3697), .ZN(n5250) );
  INV_X2 U5507 ( .A(n5247), .ZN(n3698) );
  NOR2_X2 U5508 ( .A1(n4084), .A2(n4085), .ZN(n4175) );
  INV_X2 U5510 ( .A(n5675), .ZN(n3705) );
  NOR2_X2 U5511 ( .A1(n4203), .A2(n4177), .ZN(n5672) );
  NAND3_X2 U5513 ( .A1(n3720), .A2(n3716), .A3(n3715), .ZN(\d[29] ) );
  NAND2_X2 U5514 ( .A1(n3721), .A2(n3102), .ZN(n3720) );
  OAI21_X1 U5515 ( .B1(n6360), .B2(n5677), .A(n3722), .ZN(n5673) );
  INV_X4 U5516 ( .A(n256), .ZN(n5874) );
  BUF_X4 U5517 ( .A(n3726), .Z(n3724) );
  NAND3_X2 U5518 ( .A1(n3726), .A2(n5163), .A3(n5376), .ZN(n5310) );
  XNOR2_X1 U5519 ( .A(n6016), .B(n3724), .ZN(n6018) );
  NOR2_X2 U5521 ( .A1(n2695), .A2(a[3]), .ZN(n4587) );
  NAND2_X2 U5522 ( .A1(n4328), .A2(n4329), .ZN(n4332) );
  NOR2_X2 U5523 ( .A1(n3735), .A2(n3734), .ZN(n4878) );
  AOI21_X2 U5524 ( .B1(n4813), .B2(n2734), .A(n5190), .ZN(n3734) );
  NOR2_X2 U5525 ( .A1(n4814), .A2(n4815), .ZN(n3735) );
  NOR2_X1 U5526 ( .A1(n4453), .A2(n2919), .ZN(n3737) );
  AOI21_X2 U5527 ( .B1(n342), .B2(n2907), .A(n3738), .ZN(n4487) );
  NAND2_X2 U5529 ( .A1(n3741), .A2(n4320), .ZN(n3740) );
  OAI21_X2 U5531 ( .B1(n3750), .B2(n3749), .A(n3748), .ZN(n5087) );
  INV_X2 U5532 ( .A(n3751), .ZN(n3750) );
  NAND2_X2 U5533 ( .A1(n3754), .A2(n2842), .ZN(n3753) );
  NAND2_X2 U5534 ( .A1(n5874), .A2(n5588), .ZN(n5594) );
  AOI21_X2 U5535 ( .B1(n3460), .B2(n6464), .A(n2970), .ZN(n5797) );
  AOI21_X2 U5536 ( .B1(n5785), .B2(n5784), .A(n5792), .ZN(n5786) );
  AOI22_X1 U5537 ( .A1(n4810), .A2(b[8]), .B1(n3342), .B2(n4746), .ZN(n3917)
         );
  INV_X8 U5538 ( .A(n5180), .ZN(n5266) );
  NAND2_X4 U5539 ( .A1(n5787), .A2(n5786), .ZN(n5832) );
  NAND3_X2 U5540 ( .A1(n3460), .A2(n6464), .A3(n5785), .ZN(n5787) );
  NOR2_X1 U5541 ( .A1(n4979), .A2(n4980), .ZN(n4981) );
  INV_X1 U5542 ( .A(n4883), .ZN(n4779) );
  NAND2_X1 U5543 ( .A1(n4882), .A2(n4883), .ZN(n4780) );
  NAND2_X1 U5546 ( .A1(n6011), .A2(n679), .ZN(n6012) );
  NOR2_X1 U5548 ( .A1(n5973), .A2(n2878), .ZN(n5974) );
  NAND3_X1 U5549 ( .A1(n3157), .A2(n5964), .A3(n2878), .ZN(n5965) );
  NAND2_X1 U5550 ( .A1(n5606), .A2(n2878), .ZN(n5607) );
  NAND2_X1 U5551 ( .A1(n3161), .A2(n3438), .ZN(n5001) );
  AOI22_X1 U5552 ( .A1(n4774), .A2(b[4]), .B1(n4598), .B2(n699), .ZN(n3922) );
  AND2_X4 U5553 ( .A1(n5473), .A2(n3538), .ZN(n3756) );
  XOR2_X2 U5554 ( .A(a[1]), .B(b[23]), .Z(n3757) );
  INV_X1 U5555 ( .A(n4551), .ZN(n4665) );
  XOR2_X2 U5556 ( .A(a[7]), .B(b[19]), .Z(n3763) );
  XOR2_X2 U5557 ( .A(a[13]), .B(b[11]), .Z(n3765) );
  OR4_X1 U5558 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), .ZN(n3768) );
  XNOR2_X1 U5559 ( .A(b[9]), .B(a[9]), .ZN(n3915) );
  INV_X1 U5560 ( .A(n4725), .ZN(n4679) );
  XOR2_X2 U5561 ( .A(b[7]), .B(a[23]), .Z(n4790) );
  AOI21_X1 U5562 ( .B1(n5894), .B2(n2699), .A(b[7]), .ZN(n4831) );
  XNOR2_X1 U5563 ( .A(b[19]), .B(a[19]), .ZN(n5267) );
  XNOR2_X1 U5564 ( .A(a[9]), .B(b[6]), .ZN(n3815) );
  NOR2_X1 U5565 ( .A1(b[6]), .A2(n6326), .ZN(n4499) );
  INV_X1 U5566 ( .A(n4446), .ZN(n4345) );
  INV_X1 U5567 ( .A(n4449), .ZN(n4439) );
  NAND2_X1 U5568 ( .A1(n5940), .A2(n5942), .ZN(n5912) );
  XNOR2_X1 U5569 ( .A(a[13]), .B(b[1]), .ZN(n3788) );
  INV_X1 U5570 ( .A(n5122), .ZN(n5124) );
  INV_X1 U5571 ( .A(n5272), .ZN(n5270) );
  OAI21_X1 U5572 ( .B1(n5553), .B2(n5506), .A(n5507), .ZN(n5464) );
  OAI21_X1 U5573 ( .B1(n5952), .B2(b[20]), .A(b[21]), .ZN(n5953) );
  INV_X1 U5574 ( .A(n2756), .ZN(n5157) );
  INV_X1 U5576 ( .A(n69), .ZN(n5688) );
  INV_X1 U5578 ( .A(n6117), .ZN(n6114) );
  OAI21_X1 U5579 ( .B1(n6661), .B2(n2705), .A(n5605), .ZN(n5601) );
  AOI22_X1 U5580 ( .A1(a[0]), .A2(n4128), .B1(n4219), .B2(n6569), .ZN(n5644)
         );
  AOI22_X1 U5582 ( .A1(n5856), .A2(n5924), .B1(n5855), .B2(n5854), .ZN(n5857)
         );
  NAND2_X1 U5583 ( .A1(n5980), .A2(n2878), .ZN(n5978) );
  NAND2_X1 U5586 ( .A1(n5778), .A2(n5777), .ZN(n5779) );
  INV_X8 U5593 ( .A(b[1]), .ZN(n4544) );
  NAND2_X2 U5594 ( .A1(n3952), .A2(a[15]), .ZN(n5445) );
  AOI21_X2 U5595 ( .B1(b[1]), .B2(b[0]), .A(n5445), .ZN(n3780) );
  MUX2_X2 U5596 ( .A(n1012), .B(n4405), .S(b[11]), .Z(n3784) );
  NAND2_X2 U5598 ( .A1(n2985), .A2(n3782), .ZN(n3783) );
  NOR2_X4 U5599 ( .A1(a[4]), .A2(a[3]), .ZN(n4092) );
  NAND2_X4 U5600 ( .A1(n4092), .A2(a[5]), .ZN(n4600) );
  INV_X8 U5601 ( .A(n4823), .ZN(n4601) );
  NAND2_X2 U5602 ( .A1(n3787), .A2(n3786), .ZN(n3813) );
  NAND2_X2 U5605 ( .A1(n953), .A2(n3791), .ZN(n5272) );
  NAND2_X4 U5606 ( .A1(n3793), .A2(n3792), .ZN(n4365) );
  NAND2_X2 U5607 ( .A1(n5272), .A2(n3794), .ZN(n3824) );
  NAND2_X2 U5608 ( .A1(n3799), .A2(n3798), .ZN(n4004) );
  AOI22_X2 U5610 ( .A1(n4405), .A2(b[10]), .B1(n4942), .B2(n1012), .ZN(n3808)
         );
  XNOR2_X2 U5611 ( .A(a[3]), .B(b[11]), .ZN(n3806) );
  OAI21_X2 U5612 ( .B1(n4000), .B2(n3811), .A(n3810), .ZN(n3812) );
  INV_X8 U5614 ( .A(b[14]), .ZN(n5293) );
  XOR2_X2 U5615 ( .A(a[1]), .B(b[14]), .Z(n3818) );
  AOI22_X2 U5616 ( .A1(a[0]), .A2(n3818), .B1(n4219), .B2(n4614), .ZN(n3819)
         );
  NAND2_X2 U5617 ( .A1(n3820), .A2(n3819), .ZN(n3857) );
  NAND2_X2 U5618 ( .A1(n4236), .A2(b[8]), .ZN(n3822) );
  NAND2_X4 U5620 ( .A1(a[10]), .A2(a[9]), .ZN(n5101) );
  XOR2_X2 U5623 ( .A(a[9]), .B(b[4]), .Z(n3829) );
  XOR2_X2 U5624 ( .A(a[7]), .B(b[6]), .Z(n3834) );
  XOR2_X2 U5626 ( .A(b[12]), .B(a[1]), .Z(n3839) );
  AOI22_X2 U5627 ( .A1(a[0]), .A2(n3839), .B1(n4219), .B2(n981), .ZN(n4271) );
  NOR2_X2 U5630 ( .A1(n4746), .A2(b[6]), .ZN(n3848) );
  XNOR2_X2 U5631 ( .A(b[15]), .B(a[1]), .ZN(n3850) );
  OAI22_X2 U5632 ( .A1(n3850), .A2(n4490), .B1(b[14]), .B2(n471), .ZN(n3851)
         );
  OAI21_X2 U5635 ( .B1(n3858), .B2(n3859), .A(n3857), .ZN(n3899) );
  NAND3_X2 U5637 ( .A1(n4689), .A2(a[9]), .A3(n4389), .ZN(n4609) );
  XOR2_X2 U5639 ( .A(b[16]), .B(a[1]), .Z(n3869) );
  XNOR2_X2 U5640 ( .A(a[11]), .B(b[6]), .ZN(n3871) );
  NOR2_X2 U5641 ( .A1(n4614), .A2(a[3]), .ZN(n3874) );
  NOR2_X2 U5642 ( .A1(n4492), .A2(b[13]), .ZN(n3873) );
  AOI22_X2 U5643 ( .A1(n3875), .A2(n3874), .B1(n3873), .B2(n1358), .ZN(n3876)
         );
  XNOR2_X2 U5644 ( .A(a[7]), .B(b[10]), .ZN(n3882) );
  NOR2_X2 U5645 ( .A1(n6221), .A2(a[7]), .ZN(n3879) );
  NAND2_X4 U5646 ( .A1(a[5]), .A2(a[6]), .ZN(n4948) );
  AOI21_X2 U5647 ( .B1(n3892), .B2(n3893), .A(n3891), .ZN(n3929) );
  XNOR2_X2 U5648 ( .A(a[7]), .B(b[11]), .ZN(n3962) );
  XNOR2_X2 U5649 ( .A(a[5]), .B(b[13]), .ZN(n3905) );
  XOR2_X2 U5650 ( .A(a[17]), .B(b[1]), .Z(n3906) );
  XOR2_X2 U5651 ( .A(b[17]), .B(a[1]), .Z(n3918) );
  AOI22_X2 U5652 ( .A1(a[0]), .A2(n3918), .B1(n3020), .B2(n4219), .ZN(n3943)
         );
  INV_X4 U5654 ( .A(b[4]), .ZN(n4598) );
  NOR2_X2 U5657 ( .A1(n762), .A2(n3932), .ZN(n3935) );
  NAND2_X2 U5658 ( .A1(n3932), .A2(n762), .ZN(n3934) );
  XOR2_X2 U5661 ( .A(a[15]), .B(b[4]), .Z(n3956) );
  NAND2_X2 U5662 ( .A1(n3951), .A2(b[3]), .ZN(n3953) );
  OAI22_X2 U5663 ( .A1(a[9]), .A2(n4942), .B1(n3058), .B2(b[10]), .ZN(n3960)
         );
  XOR2_X2 U5664 ( .A(a[7]), .B(b[12]), .Z(n4017) );
  XNOR2_X2 U5666 ( .A(b[18]), .B(a[1]), .ZN(n3969) );
  MUX2_X2 U5667 ( .A(n217), .B(n441), .S(b[7]), .Z(n4018) );
  XOR2_X2 U5668 ( .A(b[8]), .B(a[11]), .Z(n3970) );
  NAND2_X2 U5669 ( .A1(n2326), .A2(n3970), .ZN(n4378) );
  NOR2_X2 U5670 ( .A1(n4018), .A2(n3971), .ZN(n3972) );
  XNOR2_X2 U5671 ( .A(n3973), .B(n3972), .ZN(n3978) );
  NOR2_X2 U5672 ( .A1(n3978), .A2(n3977), .ZN(n4077) );
  INV_X4 U5675 ( .A(n4238), .ZN(n4216) );
  MUX2_X2 U5677 ( .A(n1012), .B(n4405), .S(b[9]), .Z(n3989) );
  NAND2_X2 U5679 ( .A1(a[11]), .A2(n468), .ZN(n5247) );
  NOR2_X2 U5680 ( .A1(n3992), .A2(n5247), .ZN(n4235) );
  XNOR2_X2 U5682 ( .A(b[11]), .B(a[1]), .ZN(n3995) );
  OAI21_X2 U5683 ( .B1(n3995), .B2(n4490), .A(n3994), .ZN(n3996) );
  MUX2_X2 U5684 ( .A(n6456), .B(n4601), .S(b[6]), .Z(n4245) );
  NOR2_X2 U5687 ( .A1(n4011), .A2(a[13]), .ZN(n4014) );
  XOR2_X2 U5688 ( .A(a[7]), .B(b[13]), .Z(n4016) );
  NOR3_X2 U5689 ( .A1(b[16]), .A2(a[1]), .A3(a[2]), .ZN(n4022) );
  OAI22_X2 U5690 ( .A1(n4023), .A2(a[3]), .B1(n4022), .B2(n4492), .ZN(n4024)
         );
  AOI21_X2 U5691 ( .B1(b[0]), .B2(n4030), .A(n5522), .ZN(n4031) );
  NAND2_X2 U5692 ( .A1(n1049), .A2(n1057), .ZN(n4033) );
  NOR2_X2 U5693 ( .A1(n4035), .A2(n4036), .ZN(n4037) );
  INV_X4 U5694 ( .A(n4039), .ZN(n4043) );
  AOI21_X2 U5695 ( .B1(n4043), .B2(n4042), .A(n4041), .ZN(n4376) );
  MUX2_X2 U5696 ( .A(n1354), .B(n512), .S(n4942), .Z(n4047) );
  XNOR2_X2 U5697 ( .A(a[17]), .B(b[3]), .ZN(n4049) );
  XNOR2_X2 U5698 ( .A(a[15]), .B(b[5]), .ZN(n4052) );
  OAI211_X1 U5699 ( .C1(n4065), .C2(n4064), .A(n4063), .B(n4062), .ZN(n4066)
         );
  NAND2_X2 U5700 ( .A1(n4066), .A2(n4067), .ZN(n4068) );
  NAND2_X2 U5701 ( .A1(n424), .A2(n4099), .ZN(n4088) );
  XOR2_X2 U5704 ( .A(a[3]), .B(b[4]), .Z(n4093) );
  NAND2_X2 U5705 ( .A1(n2985), .A2(n4093), .ZN(n4094) );
  MUX2_X2 U5709 ( .A(n1012), .B(n4405), .S(b[2]), .Z(n4109) );
  NAND2_X2 U5710 ( .A1(n4113), .A2(n4112), .ZN(n5662) );
  XNOR2_X2 U5711 ( .A(a[1]), .B(b[4]), .ZN(n4118) );
  MUX2_X2 U5712 ( .A(n1012), .B(n4405), .S(b[1]), .Z(n4121) );
  MUX2_X2 U5713 ( .A(n4239), .B(n4238), .S(b[2]), .Z(n4122) );
  NAND2_X2 U5715 ( .A1(a[1]), .A2(n4544), .ZN(n4125) );
  NAND2_X2 U5716 ( .A1(n4127), .A2(n4126), .ZN(n5646) );
  XOR2_X2 U5717 ( .A(b[2]), .B(a[1]), .Z(n4128) );
  NOR2_X2 U5718 ( .A1(n5646), .A2(n5644), .ZN(n6097) );
  MUX2_X2 U5719 ( .A(n1012), .B(n4405), .S(b[0]), .Z(n4130) );
  OAI21_X2 U5720 ( .B1(n4132), .B2(n4490), .A(n4131), .ZN(n4136) );
  NAND2_X2 U5721 ( .A1(n4135), .A2(n4136), .ZN(n5648) );
  NOR2_X2 U5722 ( .A1(n5652), .A2(n5648), .ZN(n5655) );
  NOR2_X2 U5723 ( .A1(n5647), .A2(n5655), .ZN(n4147) );
  NAND2_X2 U5724 ( .A1(n4134), .A2(n6096), .ZN(n5650) );
  INV_X2 U5726 ( .A(n4148), .ZN(n4146) );
  INV_X4 U5728 ( .A(n4152), .ZN(n5664) );
  AOI21_X2 U5729 ( .B1(n5667), .B2(n5664), .A(n4153), .ZN(n4155) );
  NOR2_X2 U5730 ( .A1(n5667), .A2(n5664), .ZN(n4154) );
  MUX2_X2 U5731 ( .A(n1012), .B(n4405), .S(b[5]), .Z(n4157) );
  XOR2_X2 U5732 ( .A(b[8]), .B(a[1]), .Z(n4159) );
  MUX2_X2 U5735 ( .A(n1012), .B(n4405), .S(b[6]), .Z(n4178) );
  INV_X4 U5738 ( .A(n4181), .ZN(n4182) );
  XOR2_X2 U5739 ( .A(b[9]), .B(a[1]), .Z(n4188) );
  XOR2_X2 U5740 ( .A(a[7]), .B(b[4]), .Z(n4207) );
  XOR2_X2 U5741 ( .A(a[9]), .B(b[2]), .Z(n4210) );
  MUX2_X2 U5742 ( .A(n1012), .B(n4405), .S(b[7]), .Z(n4218) );
  OAI21_X2 U5743 ( .B1(n4221), .B2(n4490), .A(n4220), .ZN(n4222) );
  NAND2_X2 U5744 ( .A1(n4223), .A2(n4222), .ZN(n4258) );
  NOR2_X2 U5745 ( .A1(n4223), .A2(n4222), .ZN(n4256) );
  MUX2_X2 U5746 ( .A(n4506), .B(n6155), .S(n3870), .Z(n4225) );
  MUX2_X2 U5747 ( .A(n1012), .B(n4405), .S(b[8]), .Z(n4237) );
  MUX2_X2 U5748 ( .A(n4239), .B(n4238), .S(b[9]), .Z(n4240) );
  NOR2_X2 U5749 ( .A1(n4241), .A2(n4240), .ZN(n4242) );
  MUX2_X2 U5750 ( .A(n1354), .B(n4795), .S(n6569), .Z(n4251) );
  OAI22_X2 U5751 ( .A1(n4252), .A2(n4251), .B1(n3035), .B2(n3037), .ZN(n4253)
         );
  AOI21_X2 U5752 ( .B1(n4257), .B2(n4258), .A(n4256), .ZN(n4288) );
  AOI22_X2 U5753 ( .A1(n4265), .A2(n4264), .B1(n4263), .B2(n4262), .ZN(n4266)
         );
  NAND2_X2 U5754 ( .A1(n1688), .A2(n4269), .ZN(n4270) );
  XNOR2_X2 U5756 ( .A(n4286), .B(n1097), .ZN(n4290) );
  INV_X2 U5757 ( .A(n1320), .ZN(n4297) );
  NOR2_X2 U5758 ( .A1(n4311), .A2(n4310), .ZN(n5704) );
  INV_X4 U5759 ( .A(n6029), .ZN(n6026) );
  XOR2_X2 U5764 ( .A(a[7]), .B(b[14]), .Z(n4334) );
  XNOR2_X2 U5766 ( .A(a[11]), .B(b[10]), .ZN(n4342) );
  XOR2_X2 U5767 ( .A(a[9]), .B(b[13]), .Z(n4346) );
  NAND2_X2 U5768 ( .A1(b[2]), .A2(n4483), .ZN(n4351) );
  XOR2_X2 U5772 ( .A(b[20]), .B(a[1]), .Z(n4361) );
  OAI22_X2 U5774 ( .A1(n4365), .A2(n4364), .B1(n4363), .B2(n4362), .ZN(n4367)
         );
  NAND2_X2 U5777 ( .A1(n4381), .A2(n4380), .ZN(n4387) );
  AOI21_X2 U5778 ( .B1(n4614), .B2(a[8]), .A(n4689), .ZN(n4391) );
  NOR2_X2 U5779 ( .A1(n4389), .A2(a[7]), .ZN(n4390) );
  OAI22_X2 U5780 ( .A1(n4391), .A2(n4390), .B1(n4998), .B2(n3638), .ZN(n4396)
         );
  NOR2_X2 U5781 ( .A1(a[9]), .A2(b[14]), .ZN(n4392) );
  NAND2_X2 U5782 ( .A1(b[14]), .A2(a[9]), .ZN(n4393) );
  NAND2_X2 U5783 ( .A1(n4394), .A2(n4393), .ZN(n4395) );
  XOR2_X2 U5784 ( .A(a[7]), .B(b[16]), .Z(n4398) );
  XOR2_X2 U5785 ( .A(a[21]), .B(b[2]), .Z(n4399) );
  BUF_X4 U5786 ( .A(n5180), .Z(n4995) );
  XNOR2_X2 U5787 ( .A(a[19]), .B(b[4]), .ZN(n4400) );
  XOR2_X2 U5789 ( .A(a[13]), .B(b[10]), .Z(n4409) );
  XNOR2_X2 U5790 ( .A(a[17]), .B(b[4]), .ZN(n4419) );
  NAND2_X2 U5793 ( .A1(a[19]), .A2(n4027), .ZN(n4425) );
  OAI22_X2 U5794 ( .A1(n4426), .A2(n4425), .B1(n4424), .B2(n4423), .ZN(n4427)
         );
  XOR2_X2 U5795 ( .A(a[13]), .B(b[9]), .Z(n4431) );
  INV_X4 U5798 ( .A(n5473), .ZN(n5526) );
  INV_X4 U5800 ( .A(n4438), .ZN(n4450) );
  OAI22_X2 U5801 ( .A1(n4441), .A2(n4440), .B1(n4450), .B2(n4439), .ZN(n4522)
         );
  XOR2_X2 U5802 ( .A(a[7]), .B(b[17]), .Z(n4482) );
  NAND3_X2 U5803 ( .A1(n4493), .A2(n1012), .A3(n4697), .ZN(n4495) );
  XNOR2_X2 U5806 ( .A(b[16]), .B(a[9]), .ZN(n4532) );
  NAND2_X2 U5809 ( .A1(a[6]), .A2(b[17]), .ZN(n4535) );
  XNOR2_X2 U5810 ( .A(a[5]), .B(b[20]), .ZN(n4540) );
  XNOR2_X2 U5811 ( .A(a[17]), .B(b[8]), .ZN(n4541) );
  OAI21_X2 U5812 ( .B1(a[23]), .B2(b[2]), .A(n4724), .ZN(n4604) );
  NOR2_X2 U5813 ( .A1(n5266), .A2(b[5]), .ZN(n4547) );
  XNOR2_X2 U5814 ( .A(a[21]), .B(b[4]), .ZN(n4548) );
  AOI21_X2 U5816 ( .B1(n5947), .B2(n4561), .A(n4560), .ZN(n4613) );
  NAND2_X2 U5818 ( .A1(b[1]), .A2(a[23]), .ZN(n4661) );
  XNOR2_X2 U5820 ( .A(a[15]), .B(b[11]), .ZN(n4595) );
  XOR2_X2 U5821 ( .A(b[5]), .B(a[21]), .Z(n4599) );
  XNOR2_X2 U5822 ( .A(a[5]), .B(b[21]), .ZN(n4602) );
  AOI22_X2 U5823 ( .A1(b[16]), .A2(n4610), .B1(n4609), .B2(n3020), .ZN(n4611)
         );
  MUX2_X2 U5824 ( .A(n5110), .B(n5109), .S(n5277), .Z(n4615) );
  NAND2_X2 U5825 ( .A1(n4621), .A2(n4622), .ZN(n4625) );
  AOI21_X2 U5828 ( .B1(n4660), .B2(a[1]), .A(n4659), .ZN(n4662) );
  MUX2_X2 U5829 ( .A(n3161), .B(n558), .S(b[13]), .Z(n4664) );
  NAND2_X2 U5830 ( .A1(n635), .A2(b[23]), .ZN(n4726) );
  NAND2_X2 U5831 ( .A1(n4678), .A2(b[23]), .ZN(n4725) );
  NOR3_X2 U5832 ( .A1(n4681), .A2(n4680), .A3(n4679), .ZN(n4682) );
  NAND2_X2 U5834 ( .A1(n4821), .A2(n3438), .ZN(n4690) );
  NOR2_X2 U5835 ( .A1(b[18]), .A2(a[9]), .ZN(n4695) );
  XOR2_X2 U5836 ( .A(a[23]), .B(b[4]), .Z(n4844) );
  OAI21_X2 U5838 ( .B1(a[3]), .B2(b[22]), .A(a[5]), .ZN(n4699) );
  AOI21_X2 U5839 ( .B1(n733), .B2(n4700), .A(n4699), .ZN(n4702) );
  XNOR2_X2 U5841 ( .A(a[11]), .B(b[16]), .ZN(n4706) );
  NAND2_X2 U5842 ( .A1(n4719), .A2(n4720), .ZN(n4722) );
  NAND3_X2 U5845 ( .A1(n4725), .A2(n4835), .A3(n6406), .ZN(n4727) );
  NAND3_X2 U5846 ( .A1(n4727), .A2(n1062), .A3(n4726), .ZN(n4728) );
  XOR2_X2 U5847 ( .A(a[15]), .B(b[13]), .Z(n4743) );
  XOR2_X2 U5848 ( .A(a[17]), .B(b[11]), .Z(n4745) );
  NOR2_X2 U5850 ( .A1(n5952), .A2(b[3]), .ZN(n4753) );
  XNOR2_X2 U5852 ( .A(a[13]), .B(b[15]), .ZN(n4755) );
  MUX2_X2 U5854 ( .A(n217), .B(n2675), .S(b[18]), .Z(n4773) );
  NAND2_X2 U5855 ( .A1(a[23]), .A2(b[4]), .ZN(n4873) );
  OAI21_X2 U5856 ( .B1(b[5]), .B2(b[4]), .A(a[23]), .ZN(n4784) );
  XNOR2_X2 U5857 ( .A(a[7]), .B(b[23]), .ZN(n4777) );
  XNOR2_X2 U5858 ( .A(a[15]), .B(b[15]), .ZN(n4788) );
  NAND2_X2 U5859 ( .A1(n4790), .A2(n5010), .ZN(n4841) );
  NAND2_X2 U5860 ( .A1(n4792), .A2(n2392), .ZN(n4953) );
  XOR2_X2 U5861 ( .A(a[9]), .B(b[22]), .Z(n4934) );
  NOR2_X2 U5863 ( .A1(n2549), .A2(n4806), .ZN(n4809) );
  XOR2_X2 U5864 ( .A(b[20]), .B(a[9]), .Z(n4811) );
  XOR2_X2 U5865 ( .A(a[7]), .B(b[22]), .Z(n4820) );
  INV_X1 U5866 ( .A(n6182), .ZN(n4818) );
  OAI22_X2 U5868 ( .A1(n4818), .A2(n4817), .B1(n4816), .B2(n4948), .ZN(n4819)
         );
  NOR2_X2 U5869 ( .A1(n4821), .A2(a[3]), .ZN(n4822) );
  XNOR2_X2 U5873 ( .A(b[8]), .B(a[21]), .ZN(n4830) );
  XNOR2_X2 U5874 ( .A(a[13]), .B(b[16]), .ZN(n4848) );
  NAND2_X2 U5875 ( .A1(n1147), .A2(b[15]), .ZN(n4850) );
  NAND2_X2 U5876 ( .A1(n4850), .A2(n4849), .ZN(n4860) );
  OAI22_X2 U5877 ( .A1(b[13]), .A2(n5076), .B1(n5077), .B2(n4614), .ZN(n4854)
         );
  NOR2_X2 U5878 ( .A1(n4852), .A2(n4851), .ZN(n4866) );
  NAND2_X2 U5880 ( .A1(n6458), .A2(n4860), .ZN(n4855) );
  XNOR2_X2 U5882 ( .A(b[8]), .B(a[23]), .ZN(n4889) );
  NOR2_X2 U5883 ( .A1(n4898), .A2(n4897), .ZN(n4926) );
  MUX2_X2 U5888 ( .A(n5074), .B(n441), .S(b[20]), .Z(n4929) );
  XOR2_X2 U5889 ( .A(a[9]), .B(b[23]), .Z(n4932) );
  XOR2_X2 U5890 ( .A(b[19]), .B(a[13]), .Z(n4941) );
  XNOR2_X2 U5891 ( .A(a[19]), .B(b[13]), .ZN(n4943) );
  NAND2_X2 U5892 ( .A1(n4944), .A2(n946), .ZN(n5016) );
  XNOR2_X2 U5893 ( .A(b[9]), .B(a[23]), .ZN(n4945) );
  XOR2_X2 U5895 ( .A(a[17]), .B(b[15]), .Z(n4949) );
  INV_X4 U5896 ( .A(n4961), .ZN(n4964) );
  XNOR2_X2 U5898 ( .A(a[17]), .B(b[16]), .ZN(n4988) );
  NAND2_X2 U5900 ( .A1(a[19]), .A2(a[20]), .ZN(n4990) );
  OAI22_X2 U5901 ( .A1(n3762), .A2(n4992), .B1(n4991), .B2(n4990), .ZN(n4993)
         );
  XOR2_X2 U5902 ( .A(a[19]), .B(b[14]), .Z(n4996) );
  NAND2_X2 U5903 ( .A1(a[23]), .A2(b[8]), .ZN(n5044) );
  XNOR2_X2 U5905 ( .A(a[15]), .B(b[18]), .ZN(n5003) );
  NAND2_X2 U5906 ( .A1(n6221), .A2(a[23]), .ZN(n5007) );
  NAND2_X2 U5907 ( .A1(n5952), .A2(b[9]), .ZN(n5006) );
  INV_X4 U5911 ( .A(n5042), .ZN(n5043) );
  NAND2_X2 U5912 ( .A1(n5043), .A2(n3632), .ZN(n5046) );
  MUX2_X2 U5913 ( .A(n699), .B(n4774), .S(b[20]), .Z(n5049) );
  MUX2_X2 U5914 ( .A(n1318), .B(n5900), .S(b[10]), .Z(n5057) );
  OAI22_X2 U5915 ( .A1(n5068), .A2(n5067), .B1(n5066), .B2(n6153), .ZN(n5133)
         );
  NOR2_X2 U5916 ( .A1(n5071), .A2(n610), .ZN(n5466) );
  MUX2_X2 U5917 ( .A(n5074), .B(n440), .S(b[22]), .Z(n5075) );
  OAI21_X2 U5919 ( .B1(b[8]), .B2(b[9]), .A(a[23]), .ZN(n5151) );
  INV_X4 U5920 ( .A(n5087), .ZN(n5088) );
  INV_X4 U5922 ( .A(n5622), .ZN(n5376) );
  NAND3_X2 U5923 ( .A1(b[23]), .A2(a[10]), .A3(n5100), .ZN(n5103) );
  NAND2_X2 U5925 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  NAND2_X2 U5927 ( .A1(n5106), .A2(b[22]), .ZN(n5107) );
  MUX2_X2 U5929 ( .A(n5110), .B(n5109), .S(n5951), .Z(n5165) );
  NOR2_X2 U5930 ( .A1(n5117), .A2(n4046), .ZN(n5120) );
  OAI22_X2 U5932 ( .A1(n5125), .A2(n5124), .B1(n5123), .B2(n1805), .ZN(n5128)
         );
  XOR2_X2 U5935 ( .A(a[21]), .B(b[14]), .Z(n5137) );
  MUX2_X2 U5936 ( .A(n6035), .B(n5899), .S(b[12]), .Z(n5141) );
  MUX2_X2 U5937 ( .A(n5947), .B(n5900), .S(b[11]), .Z(n5140) );
  XNOR2_X2 U5939 ( .A(a[17]), .B(b[18]), .ZN(n5148) );
  XNOR2_X2 U5940 ( .A(n5186), .B(n5187), .ZN(n5152) );
  OAI21_X2 U5943 ( .B1(n833), .B2(n5159), .A(n5158), .ZN(n5315) );
  AOI21_X2 U5944 ( .B1(n5620), .B2(n5376), .A(n5160), .ZN(n5602) );
  NAND2_X2 U5945 ( .A1(b[11]), .A2(b[10]), .ZN(n5241) );
  OAI21_X2 U5946 ( .B1(b[11]), .B2(b[10]), .A(a[23]), .ZN(n5240) );
  XOR2_X2 U5947 ( .A(b[17]), .B(a[19]), .Z(n5178) );
  XOR2_X2 U5948 ( .A(a[13]), .B(b[23]), .Z(n5184) );
  NOR2_X2 U5949 ( .A1(n5192), .A2(n5191), .ZN(n5229) );
  XOR2_X2 U5950 ( .A(b[15]), .B(a[21]), .Z(n5193) );
  MUX2_X2 U5951 ( .A(n5077), .B(n5076), .S(n5471), .Z(n5199) );
  NOR2_X1 U5952 ( .A1(n5079), .A2(n5196), .ZN(n5198) );
  NOR2_X2 U5953 ( .A1(n5199), .A2(n5198), .ZN(n5228) );
  OAI21_X2 U5954 ( .B1(n5211), .B2(n5210), .A(n5209), .ZN(n5215) );
  NAND2_X2 U5956 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  NAND2_X2 U5957 ( .A1(n5225), .A2(n6674), .ZN(n5230) );
  AOI22_X2 U5958 ( .A1(n5230), .A2(n5229), .B1(n5228), .B2(n5227), .ZN(n5289)
         );
  XNOR2_X2 U5960 ( .A(a[17]), .B(b[20]), .ZN(n5233) );
  MUX2_X2 U5961 ( .A(n4995), .B(n465), .S(b[17]), .Z(n5236) );
  NAND2_X2 U5962 ( .A1(n5237), .A2(n5236), .ZN(n5285) );
  MUX2_X2 U5963 ( .A(n1761), .B(n5136), .S(b[15]), .Z(n5245) );
  XOR2_X2 U5964 ( .A(b[16]), .B(a[21]), .Z(n5243) );
  NAND2_X2 U5965 ( .A1(n3334), .A2(n5243), .ZN(n5244) );
  NAND2_X2 U5966 ( .A1(n5245), .A2(n5244), .ZN(n5298) );
  AOI22_X2 U5967 ( .A1(n5250), .A2(n5249), .B1(n888), .B2(n3698), .ZN(n5297)
         );
  OAI21_X2 U5969 ( .B1(n5256), .B2(n6424), .A(n5254), .ZN(n5264) );
  NOR2_X2 U5970 ( .A1(n716), .A2(n637), .ZN(n5628) );
  NAND2_X2 U5971 ( .A1(n5272), .A2(n5273), .ZN(n5349) );
  MUX2_X2 U5972 ( .A(n5077), .B(n5076), .S(n566), .Z(n5274) );
  MUX2_X2 U5973 ( .A(n1194), .B(n1193), .S(n5471), .Z(n5275) );
  MUX2_X2 U5974 ( .A(n5294), .B(n5278), .S(b[13]), .Z(n5279) );
  NAND2_X2 U5975 ( .A1(n5280), .A2(n5281), .ZN(n5357) );
  NAND2_X2 U5976 ( .A1(n5357), .A2(n5356), .ZN(n5287) );
  INV_X4 U5978 ( .A(n6035), .ZN(n5476) );
  INV_X4 U5979 ( .A(n5297), .ZN(n5300) );
  NAND2_X2 U5980 ( .A1(n5300), .A2(n6154), .ZN(n5302) );
  NOR2_X2 U5981 ( .A1(n5300), .A2(n6154), .ZN(n5301) );
  NOR2_X2 U5982 ( .A1(n5319), .A2(n5318), .ZN(n5971) );
  NAND3_X2 U5984 ( .A1(n5310), .A2(n5602), .A3(n6526), .ZN(n5314) );
  INV_X4 U5985 ( .A(n5315), .ZN(n5316) );
  BUF_X4 U5986 ( .A(n6071), .Z(n5998) );
  OAI21_X2 U5987 ( .B1(n660), .B2(n5334), .A(n5333), .ZN(n5371) );
  NOR2_X1 U5988 ( .A1(n5337), .A2(b[23]), .ZN(n5338) );
  AOI21_X2 U5990 ( .B1(n5345), .B2(n5344), .A(n5343), .ZN(n5346) );
  MUX2_X2 U5992 ( .A(n6035), .B(n5899), .S(b[16]), .Z(n5359) );
  MUX2_X2 U5993 ( .A(n1318), .B(n5900), .S(b[15]), .Z(n5358) );
  NAND2_X2 U5994 ( .A1(n5364), .A2(n5363), .ZN(n5366) );
  INV_X4 U5995 ( .A(n5371), .ZN(n5372) );
  NAND2_X2 U5996 ( .A1(n3476), .A2(n5378), .ZN(n5379) );
  NAND2_X2 U5997 ( .A1(n5388), .A2(n5387), .ZN(n5392) );
  NAND2_X2 U5999 ( .A1(n5420), .A2(n5397), .ZN(n5399) );
  NAND2_X2 U6000 ( .A1(n5399), .A2(n5398), .ZN(n5403) );
  MUX2_X2 U6001 ( .A(n5948), .B(n5476), .S(n5471), .Z(n5401) );
  BUF_X4 U6002 ( .A(n4752), .Z(n6043) );
  MUX2_X2 U6003 ( .A(n6043), .B(n3142), .S(n3438), .Z(n5400) );
  NOR2_X2 U6004 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  NOR2_X2 U6005 ( .A1(n5403), .A2(n5402), .ZN(n5537) );
  NAND2_X2 U6006 ( .A1(n5403), .A2(n5402), .ZN(n5535) );
  NAND2_X2 U6007 ( .A1(n5404), .A2(n5535), .ZN(n5408) );
  MUX2_X2 U6008 ( .A(n5948), .B(n5476), .S(n3438), .Z(n5406) );
  MUX2_X2 U6009 ( .A(n6043), .B(n3142), .S(n5360), .Z(n5405) );
  NOR2_X2 U6010 ( .A1(n5406), .A2(n5405), .ZN(n5416) );
  AOI21_X2 U6011 ( .B1(n3766), .B2(n5416), .A(n5407), .ZN(n5536) );
  XOR2_X2 U6012 ( .A(n5408), .B(n5536), .Z(n5413) );
  NAND2_X2 U6013 ( .A1(a[23]), .A2(b[18]), .ZN(n5531) );
  NAND2_X2 U6014 ( .A1(n5413), .A2(n5412), .ZN(n5539) );
  NAND2_X2 U6015 ( .A1(n5414), .A2(n5539), .ZN(n5432) );
  XNOR2_X2 U6016 ( .A(n5417), .B(n5416), .ZN(n5430) );
  XNOR2_X2 U6017 ( .A(n5420), .B(n5419), .ZN(n5429) );
  NOR2_X2 U6018 ( .A1(n5430), .A2(n5429), .ZN(n5421) );
  NAND2_X2 U6019 ( .A1(n5430), .A2(n5429), .ZN(n5433) );
  AOI21_X2 U6020 ( .B1(n5434), .B2(n5435), .A(n5431), .ZN(n5540) );
  NOR2_X2 U6021 ( .A1(n5441), .A2(n5440), .ZN(n5496) );
  MUX2_X2 U6023 ( .A(n5947), .B(n5900), .S(b[16]), .Z(n5443) );
  AOI21_X2 U6024 ( .B1(n5444), .B2(n5443), .A(n5442), .ZN(n5494) );
  NAND2_X2 U6025 ( .A1(n5444), .A2(n5443), .ZN(n5446) );
  NOR2_X2 U6026 ( .A1(n5446), .A2(n5445), .ZN(n5495) );
  MUX2_X2 U6027 ( .A(n314), .B(n5454), .S(b[23]), .Z(n5456) );
  NAND2_X2 U6029 ( .A1(n5462), .A2(n5461), .ZN(n5502) );
  NOR2_X2 U6030 ( .A1(n5468), .A2(n5467), .ZN(n5500) );
  AOI21_X2 U6031 ( .B1(n5500), .B2(n5470), .A(n5469), .ZN(n5511) );
  MUX2_X2 U6032 ( .A(n5472), .B(n5897), .S(n5471), .Z(n5475) );
  MUX2_X2 U6033 ( .A(n3230), .B(n5136), .S(b[19]), .Z(n5474) );
  NAND2_X2 U6034 ( .A1(n5475), .A2(n5474), .ZN(n5510) );
  MUX2_X2 U6035 ( .A(n5948), .B(n5476), .S(n5360), .Z(n5479) );
  MUX2_X2 U6036 ( .A(n6043), .B(n3142), .S(n3217), .Z(n5478) );
  NOR2_X2 U6037 ( .A1(n5479), .A2(n5478), .ZN(n5509) );
  AOI21_X2 U6038 ( .B1(n5483), .B2(n5482), .A(n5481), .ZN(n5484) );
  NOR2_X2 U6039 ( .A1(n5495), .A2(n5494), .ZN(n5497) );
  XNOR2_X2 U6040 ( .A(n5500), .B(n5499), .ZN(n5501) );
  XNOR2_X2 U6041 ( .A(n5510), .B(n5509), .ZN(n5512) );
  XNOR2_X2 U6042 ( .A(n5512), .B(n5511), .ZN(n5513) );
  AOI21_X2 U6043 ( .B1(n5548), .B2(n5546), .A(n5515), .ZN(n5572) );
  NOR2_X2 U6044 ( .A1(n5914), .A2(n5913), .ZN(n6063) );
  MUX2_X2 U6045 ( .A(n6035), .B(n5899), .S(b[21]), .Z(n5519) );
  MUX2_X2 U6046 ( .A(n5947), .B(n5900), .S(b[20]), .Z(n5518) );
  NAND2_X2 U6047 ( .A1(n5519), .A2(n5518), .ZN(n5523) );
  NAND2_X2 U6048 ( .A1(n5521), .A2(n5520), .ZN(n5942) );
  NAND2_X2 U6050 ( .A1(n5942), .A2(n5892), .ZN(n5524) );
  XNOR2_X2 U6051 ( .A(n5893), .B(n5524), .ZN(n5534) );
  NOR2_X2 U6052 ( .A1(n5528), .A2(n5527), .ZN(n5906) );
  XNOR2_X2 U6053 ( .A(n5906), .B(n5532), .ZN(n5533) );
  OAI21_X2 U6054 ( .B1(n5541), .B2(n5540), .A(n5539), .ZN(n5544) );
  NAND2_X2 U6055 ( .A1(n5543), .A2(n5542), .ZN(n6077) );
  NAND2_X2 U6056 ( .A1(n6077), .A2(n6064), .ZN(n5575) );
  NAND2_X2 U6057 ( .A1(n6063), .A2(n5575), .ZN(n5583) );
  NOR2_X2 U6058 ( .A1(n5552), .A2(n5551), .ZN(n5554) );
  NAND2_X2 U6059 ( .A1(n5560), .A2(n5559), .ZN(n5579) );
  INV_X4 U6060 ( .A(n5875), .ZN(n5915) );
  NOR2_X2 U6061 ( .A1(n5915), .A2(n5570), .ZN(n5612) );
  NAND2_X2 U6062 ( .A1(n5569), .A2(n6072), .ZN(n5590) );
  NAND2_X2 U6064 ( .A1(n2725), .A2(n5574), .ZN(n6068) );
  INV_X4 U6065 ( .A(n6068), .ZN(n5933) );
  NOR2_X2 U6066 ( .A1(n5933), .A2(n5575), .ZN(n5582) );
  NOR2_X2 U6067 ( .A1(n5591), .A2(n6072), .ZN(n5585) );
  AOI21_X2 U6068 ( .B1(n5589), .B2(n5588), .A(n3768), .ZN(n5595) );
  INV_X1 U6069 ( .A(n5599), .ZN(n5600) );
  NAND3_X2 U6071 ( .A1(n5885), .A2(n5616), .A3(n3164), .ZN(n5614) );
  NOR2_X2 U6072 ( .A1(n5612), .A2(n5611), .ZN(n5615) );
  NAND2_X2 U6073 ( .A1(n5614), .A2(n5613), .ZN(n5619) );
  NAND2_X2 U6075 ( .A1(n5969), .A2(n5975), .ZN(n5634) );
  NAND2_X2 U6077 ( .A1(n5976), .A2(n5634), .ZN(n5638) );
  NOR2_X1 U6078 ( .A1(n1355), .A2(n259), .ZN(n5637) );
  OAI22_X2 U6079 ( .A1(n6056), .A2(n5638), .B1(n5637), .B2(n5636), .ZN(n5639)
         );
  NOR3_X2 U6080 ( .A1(n5641), .A2(n5640), .A3(n5639), .ZN(\d[36]_BAR ) );
  NOR2_X2 U6083 ( .A1(n5683), .A2(n325), .ZN(n5696) );
  NOR2_X2 U6084 ( .A1(n5684), .A2(n5696), .ZN(n5687) );
  NOR2_X2 U6085 ( .A1(n5710), .A2(n3167), .ZN(n5708) );
  NAND2_X2 U6086 ( .A1(n5715), .A2(n5714), .ZN(n5720) );
  NAND2_X4 U6087 ( .A1(n5725), .A2(n5724), .ZN(n5778) );
  NAND2_X2 U6088 ( .A1(n5726), .A2(n5778), .ZN(n5728) );
  NAND2_X2 U6091 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  NAND2_X2 U6092 ( .A1(n5738), .A2(n5739), .ZN(\d[17]_BAR ) );
  NOR2_X2 U6093 ( .A1(n5741), .A2(n5740), .ZN(n5760) );
  INV_X4 U6094 ( .A(n2970), .ZN(n5783) );
  NAND2_X2 U6095 ( .A1(n5748), .A2(n5783), .ZN(n5747) );
  NOR2_X2 U6096 ( .A1(n5744), .A2(n5743), .ZN(n5756) );
  NOR2_X2 U6097 ( .A1(n5746), .A2(n5745), .ZN(n5758) );
  NOR2_X2 U6098 ( .A1(n5749), .A2(n5748), .ZN(n5753) );
  NAND3_X2 U6099 ( .A1(n5756), .A2(n5755), .A3(n5754), .ZN(\d[19] ) );
  NAND2_X2 U6100 ( .A1(n5758), .A2(n5778), .ZN(n5759) );
  AOI21_X2 U6101 ( .B1(n5759), .B2(n5760), .A(n143), .ZN(n5762) );
  NAND2_X2 U6102 ( .A1(n5762), .A2(n5763), .ZN(n5761) );
  OAI21_X2 U6103 ( .B1(n5763), .B2(n5762), .A(n5761), .ZN(\d[18] ) );
  OAI21_X2 U6104 ( .B1(n5766), .B2(n5773), .A(n5765), .ZN(n5770) );
  XNOR2_X2 U6105 ( .A(n5770), .B(n5769), .ZN(\d[16] ) );
  BUF_X4 U6107 ( .A(n5780), .Z(n5799) );
  NOR2_X2 U6108 ( .A1(n5781), .A2(n5799), .ZN(n5791) );
  NOR2_X2 U6109 ( .A1(n5796), .A2(n5791), .ZN(n5785) );
  BUF_X4 U6110 ( .A(n5805), .Z(n5806) );
  OAI21_X2 U6111 ( .B1(n3427), .B2(n5838), .A(n6375), .ZN(n5811) );
  INV_X1 U6112 ( .A(n2681), .ZN(n5824) );
  AOI21_X2 U6113 ( .B1(n5824), .B2(n5821), .A(n5814), .ZN(n5829) );
  AOI21_X2 U6114 ( .B1(n5832), .B2(n5816), .A(n5815), .ZN(n5820) );
  AOI21_X2 U6115 ( .B1(n5832), .B2(n6453), .A(n5821), .ZN(n5826) );
  AOI21_X2 U6116 ( .B1(n5832), .B2(n5831), .A(n5830), .ZN(n5833) );
  NOR2_X2 U6119 ( .A1(n3552), .A2(n5858), .ZN(n5843) );
  INV_X1 U6120 ( .A(n5851), .ZN(n5852) );
  XNOR2_X2 U6121 ( .A(n5859), .B(n3679), .ZN(n5861) );
  NOR2_X2 U6124 ( .A1(n5933), .A2(n5914), .ZN(n5878) );
  INV_X4 U6125 ( .A(n679), .ZN(n6062) );
  NOR2_X2 U6126 ( .A1(n5878), .A2(n5913), .ZN(n5882) );
  NAND2_X2 U6127 ( .A1(n5882), .A2(n1314), .ZN(n5884) );
  NAND2_X2 U6128 ( .A1(n5877), .A2(n5878), .ZN(n5880) );
  OAI22_X2 U6129 ( .A1(n6070), .A2(n5880), .B1(n5994), .B2(n5879), .ZN(n5881)
         );
  NOR2_X2 U6130 ( .A1(n5394), .A2(n5927), .ZN(n5921) );
  MUX2_X2 U6131 ( .A(n5896), .B(n5136), .S(b[23]), .Z(n5898) );
  NAND2_X2 U6132 ( .A1(n5898), .A2(n5897), .ZN(n5958) );
  XNOR2_X2 U6133 ( .A(n5958), .B(n5957), .ZN(n5903) );
  MUX2_X2 U6134 ( .A(n195), .B(n5899), .S(b[22]), .Z(n5902) );
  MUX2_X2 U6135 ( .A(n6585), .B(n5900), .S(b[21]), .Z(n5901) );
  NAND2_X2 U6136 ( .A1(n5902), .A2(n5901), .ZN(n5956) );
  XNOR2_X2 U6137 ( .A(n5903), .B(n5956), .ZN(n5907) );
  AOI21_X2 U6138 ( .B1(n5906), .B2(n5905), .A(n5904), .ZN(n5908) );
  NAND2_X2 U6139 ( .A1(n5907), .A2(n5908), .ZN(n5939) );
  NAND2_X2 U6140 ( .A1(n5910), .A2(n5909), .ZN(n5941) );
  NAND2_X2 U6141 ( .A1(n5939), .A2(n5941), .ZN(n5911) );
  NOR2_X2 U6142 ( .A1(n5918), .A2(n5917), .ZN(n5920) );
  NOR3_X2 U6143 ( .A1(n5946), .A2(n5945), .A3(n5944), .ZN(n6112) );
  OAI22_X2 U6144 ( .A1(n195), .A2(b[23]), .B1(b[22]), .B2(n6585), .ZN(n6032)
         );
  XNOR2_X2 U6145 ( .A(n5955), .B(n5954), .ZN(n6027) );
  AOI22_X2 U6147 ( .A1(n5961), .A2(n5960), .B1(n6033), .B2(n5959), .ZN(n6030)
         );
  XNOR2_X2 U6148 ( .A(n5962), .B(n6030), .ZN(n6117) );
  NAND2_X2 U6149 ( .A1(n6058), .A2(n5964), .ZN(n5967) );
  NAND2_X2 U6151 ( .A1(n5970), .A2(n5969), .ZN(n5981) );
  NOR2_X2 U6152 ( .A1(n5981), .A2(n5977), .ZN(n5984) );
  NAND2_X2 U6153 ( .A1(n5976), .A2(n5975), .ZN(n5985) );
  NOR2_X2 U6154 ( .A1(n5985), .A2(n5983), .ZN(n5980) );
  NAND2_X2 U6155 ( .A1(n5979), .A2(n5978), .ZN(n5993) );
  NOR2_X2 U6157 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  NAND2_X2 U6158 ( .A1(n5995), .A2(n5994), .ZN(n6001) );
  NAND2_X2 U6159 ( .A1(n5996), .A2(n6001), .ZN(n6006) );
  XNOR2_X2 U6165 ( .A(n6048), .B(n6101), .ZN(n6121) );
  AOI21_X2 U6169 ( .B1(n6059), .B2(n6058), .A(n6057), .ZN(n6060) );
  NAND2_X2 U6170 ( .A1(n6060), .A2(n6061), .ZN(\d[46]_BAR ) );
  OAI211_X1 U6171 ( .C1(n6068), .C2(n6067), .A(n6066), .B(n6077), .ZN(n6069)
         );
  AOI21_X2 U6172 ( .B1(n6070), .B2(n6073), .A(n6069), .ZN(n6080) );
  AOI21_X2 U6174 ( .B1(n6166), .B2(n6080), .A(n3767), .ZN(n6082) );
  OAI21_X2 U6175 ( .B1(n496), .B2(n6083), .A(n6082), .ZN(n6091) );
  NOR2_X2 U6176 ( .A1(n61), .A2(n6085), .ZN(n6087) );
  NAND2_X2 U6177 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  INV_X2 U6178 ( .A(n6089), .ZN(n6090) );
  NOR2_X2 U6179 ( .A1(n6091), .A2(n6090), .ZN(\d[44] ) );
  XOR2_X1 U6180 ( .A(n6093), .B(n6092), .Z(n6095) );
  INV_X1 U6181 ( .A(n6099), .ZN(n6100) );
  MUX2_X2 U6182 ( .A(n6103), .B(n6102), .S(n6101), .Z(n6106) );
  NOR2_X2 U6183 ( .A1(n6110), .A2(n6115), .ZN(n6133) );
  INV_X4 U3626 ( .A(n4314), .ZN(n4007) );
  NAND2_X2 U1216 ( .A1(n295), .A2(n296), .ZN(n298) );
  AOI21_X2 U1214 ( .B1(n4231), .B2(n4232), .A(n1124), .ZN(n4260) );
  NAND3_X2 U980 ( .A1(n4937), .A2(n4938), .A3(n4939), .ZN(n209) );
  INV_X8 U4782 ( .A(n440), .ZN(n4705) );
  NOR2_X2 U4771 ( .A1(n5293), .A2(n4590), .ZN(n4591) );
  NOR2_X2 U2052 ( .A1(n5032), .A2(n3379), .ZN(n3378) );
  XNOR2_X2 U4849 ( .A(n5635), .B(n1355), .ZN(n5636) );
  INV_X4 U1302 ( .A(n5258), .ZN(n5257) );
  OAI21_X2 U3775 ( .B1(n2573), .B2(n6198), .A(n3620), .ZN(n1664) );
  NOR2_X4 U3500 ( .A1(n2489), .A2(n954), .ZN(n1391) );
  NAND2_X4 U1303 ( .A1(n5258), .A2(n6165), .ZN(n5262) );
  NAND2_X2 U2275 ( .A1(n1700), .A2(n1019), .ZN(n868) );
  INV_X2 U294 ( .A(n28), .ZN(n46) );
  NAND2_X2 U1903 ( .A1(n5293), .A2(n6457), .ZN(n3500) );
  AOI21_X2 U1589 ( .B1(n4457), .B2(n4456), .A(n4455), .ZN(n4469) );
  NOR3_X2 U157 ( .A1(n6413), .A2(n4982), .A3(n5845), .ZN(n4970) );
  NAND2_X4 U1237 ( .A1(n5262), .A2(n5261), .ZN(n5309) );
  NAND2_X2 U521 ( .A1(n1847), .A2(n2244), .ZN(n2994) );
  INV_X4 U4024 ( .A(n6155), .ZN(n3614) );
  NOR2_X4 U5337 ( .A1(n3352), .A2(n5894), .ZN(n6029) );
  INV_X4 U4517 ( .A(n139), .ZN(n4806) );
  INV_X4 U4128 ( .A(n2042), .ZN(n3256) );
  INV_X4 U2246 ( .A(n1485), .ZN(n848) );
  NAND2_X4 U37 ( .A1(n1568), .A2(n1567), .ZN(n4445) );
  INV_X4 U4986 ( .A(n3557), .ZN(n4895) );
  INV_X4 U1966 ( .A(n1468), .ZN(n662) );
  NOR2_X4 U707 ( .A1(n1940), .A2(n138), .ZN(n1468) );
  OAI21_X2 U1126 ( .B1(n4575), .B2(n4574), .A(n4573), .ZN(n4627) );
  INV_X4 U754 ( .A(n3273), .ZN(n151) );
  INV_X2 U2072 ( .A(n2930), .ZN(n737) );
  AOI21_X2 U4778 ( .B1(n5110), .B2(b[17]), .A(n2850), .ZN(n2849) );
  NAND2_X2 U2202 ( .A1(b[18]), .A2(n5041), .ZN(n2501) );
  INV_X4 U3648 ( .A(n1625), .ZN(n5053) );
  NOR2_X2 U3101 ( .A1(n3210), .A2(n1148), .ZN(n4766) );
  NAND2_X2 U2245 ( .A1(n5899), .A2(b[14]), .ZN(n3514) );
  NOR3_X4 U5420 ( .A1(n4812), .A2(a[23]), .A3(n6328), .ZN(n3512) );
  INV_X4 U2788 ( .A(n5284), .ZN(n1037) );
  AOI22_X2 U1196 ( .A1(n5525), .A2(b[17]), .B1(n3020), .B2(n5526), .ZN(n2053)
         );
  NAND2_X2 U519 ( .A1(n3079), .A2(n4627), .ZN(n85) );
  OAI21_X2 U4219 ( .B1(n6155), .B2(b[16]), .A(n2161), .ZN(n4319) );
  INV_X4 U5322 ( .A(n3858), .ZN(n3301) );
  OAI21_X2 U2271 ( .B1(n1464), .B2(n2584), .A(n4936), .ZN(n1463) );
  INV_X4 U2606 ( .A(n2584), .ZN(n1011) );
  INV_X4 U5402 ( .A(a[15]), .ZN(n3951) );
  NOR2_X2 U1487 ( .A1(n4442), .A2(n2042), .ZN(n2041) );
  NAND2_X2 U4826 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  NAND2_X2 U2095 ( .A1(n1847), .A2(n5360), .ZN(n3643) );
  XOR2_X2 U2374 ( .A(b[10]), .B(a[23]), .Z(n5009) );
  XNOR2_X2 U2375 ( .A(a[13]), .B(b[6]), .ZN(n3968) );
  INV_X4 U90 ( .A(b[18]), .ZN(n5360) );
  INV_X4 U5762 ( .A(n4329), .ZN(n4330) );
  NOR2_X4 U64 ( .A1(n6589), .A2(n4709), .ZN(n2965) );
  NAND2_X2 U2402 ( .A1(n6203), .A2(b[3]), .ZN(n4209) );
  OAI21_X2 U1946 ( .B1(n4234), .B2(n69), .A(n4233), .ZN(n5685) );
  INV_X8 U5059 ( .A(a[17]), .ZN(n2909) );
  NAND2_X4 U527 ( .A1(n2022), .A2(n2833), .ZN(n1543) );
  NAND2_X2 U2070 ( .A1(n5050), .A2(n5049), .ZN(n2759) );
  NOR2_X2 U3889 ( .A1(n1308), .A2(b[7]), .ZN(n2212) );
  NAND2_X2 U1569 ( .A1(n3629), .A2(n2757), .ZN(n1283) );
  INV_X4 U4258 ( .A(n3859), .ZN(n2210) );
  INV_X4 U3983 ( .A(n3399), .ZN(n3312) );
  INV_X8 U3761 ( .A(n4829), .ZN(n5136) );
  NOR2_X2 U1515 ( .A1(n4593), .A2(n2327), .ZN(n4594) );
  NAND3_X4 U1734 ( .A1(n1916), .A2(a[12]), .A3(a[11]), .ZN(n558) );
  NAND3_X2 U5056 ( .A1(n3476), .A2(n628), .A3(n343), .ZN(n5923) );
  NOR2_X2 U4751 ( .A1(n6185), .A2(n2380), .ZN(n4023) );
  NAND2_X2 U1317 ( .A1(n2636), .A2(n1367), .ZN(n338) );
  NOR2_X4 U4245 ( .A1(n414), .A2(n2716), .ZN(n2199) );
  NAND2_X4 U2508 ( .A1(n1539), .A2(n4086), .ZN(n4099) );
  NAND2_X2 U1287 ( .A1(n4219), .A2(n3835), .ZN(n4086) );
  NAND2_X2 U1422 ( .A1(n396), .A2(n1151), .ZN(n1150) );
  NAND2_X2 U2166 ( .A1(n184), .A2(n4239), .ZN(n1738) );
  NOR2_X4 U544 ( .A1(n4503), .A2(n3439), .ZN(n2484) );
  NOR2_X4 U565 ( .A1(n3430), .A2(n2485), .ZN(n3439) );
  NAND2_X1 U1204 ( .A1(n5053), .A2(n5054), .ZN(n1515) );
  OAI22_X2 U2334 ( .A1(n4418), .A2(n4490), .B1(b[21]), .B2(n472), .ZN(n4497)
         );
  NAND2_X4 U2278 ( .A1(n870), .A2(n5256), .ZN(n872) );
  NAND2_X2 U1342 ( .A1(n4019), .A2(n4020), .ZN(n352) );
  NOR2_X4 U5499 ( .A1(n4794), .A2(n3438), .ZN(n3685) );
  INV_X4 U3625 ( .A(n1751), .ZN(n5030) );
  AOI21_X2 U3142 ( .B1(n2066), .B2(n4885), .A(n4884), .ZN(n4918) );
  INV_X4 U1479 ( .A(n6328), .ZN(n2513) );
  INV_X4 U2633 ( .A(b[16]), .ZN(n2380) );
  AOI21_X2 U4856 ( .B1(n5882), .B2(n6070), .A(n5881), .ZN(n5883) );
  NAND2_X2 U2060 ( .A1(n5562), .A2(n5561), .ZN(n731) );
  NAND2_X2 U5520 ( .A1(n4581), .A2(n3492), .ZN(n4639) );
  NAND2_X2 U2270 ( .A1(n2586), .A2(n2585), .ZN(n3104) );
  NOR2_X2 U5482 ( .A1(b[1]), .A2(n4600), .ZN(n3665) );
  NAND2_X4 U1563 ( .A1(n466), .A2(n359), .ZN(n469) );
  NOR2_X4 U912 ( .A1(n3685), .A2(n1329), .ZN(n193) );
  NAND2_X4 U1564 ( .A1(n360), .A2(n469), .ZN(n2889) );
  NOR2_X4 U629 ( .A1(n5234), .A2(n113), .ZN(n5283) );
  NAND2_X2 U2195 ( .A1(n1880), .A2(n814), .ZN(n815) );
  AOI21_X2 U4766 ( .B1(n2249), .B2(n5076), .A(n2997), .ZN(n2996) );
  XOR2_X2 U1748 ( .A(n2695), .B(n4661), .Z(n2714) );
  OAI21_X2 U1738 ( .B1(n4462), .B2(n4469), .A(n6495), .ZN(n4471) );
  XOR2_X2 U2380 ( .A(b[20]), .B(a[11]), .Z(n2701) );
  INV_X2 U2925 ( .A(b[1]), .ZN(n3367) );
  NAND2_X2 U4862 ( .A1(b[1]), .A2(a[0]), .ZN(n5643) );
  INV_X4 U2526 ( .A(b[16]), .ZN(n3020) );
  INV_X2 U2910 ( .A(b[23]), .ZN(n3154) );
  INV_X2 U2905 ( .A(b[23]), .ZN(n1896) );
  XNOR2_X1 U2384 ( .A(b[20]), .B(a[13]), .ZN(n5002) );
  INV_X4 U102 ( .A(b[0]), .ZN(n2603) );
  XOR2_X2 U2383 ( .A(a[9]), .B(b[15]), .Z(n4481) );
  INV_X2 U2390 ( .A(b[23]), .ZN(n5221) );
  XOR2_X2 U5588 ( .A(n5643), .B(n5642), .Z(\d[1] ) );
  AND2_X2 U2424 ( .A1(n3022), .A2(b[16]), .ZN(n955) );
  NAND2_X2 U2014 ( .A1(n703), .A2(n704), .ZN(n706) );
  NOR2_X1 U4260 ( .A1(n6203), .A2(n3465), .ZN(n2213) );
  NAND2_X2 U1877 ( .A1(n624), .A2(n625), .ZN(n627) );
  AND2_X1 U2514 ( .A1(n3632), .A2(b[9]), .ZN(n5150) );
  INV_X2 U5849 ( .A(n4754), .ZN(n4751) );
  NAND2_X2 U4176 ( .A1(n2335), .A2(n3540), .ZN(n4160) );
  NOR2_X2 U1174 ( .A1(n4930), .A2(n4929), .ZN(n3269) );
  INV_X2 U4381 ( .A(n2371), .ZN(n2370) );
  AND2_X2 U1550 ( .A1(n3562), .A2(n530), .ZN(n464) );
  INV_X2 U2415 ( .A(n4789), .ZN(n4791) );
  INV_X2 U1382 ( .A(n4452), .ZN(n379) );
  INV_X2 U254 ( .A(n2868), .ZN(n19) );
  NAND2_X2 U5466 ( .A1(n3624), .A2(n3623), .ZN(n3622) );
  INV_X2 U5770 ( .A(n2906), .ZN(n4352) );
  INV_X2 U499 ( .A(n4510), .ZN(n4508) );
  NOR2_X2 U1116 ( .A1(n5005), .A2(n5004), .ZN(n5054) );
  NAND2_X2 U53 ( .A1(n3805), .A2(n3804), .ZN(n4000) );
  OR2_X2 U2427 ( .A1(n4272), .A2(n3425), .ZN(n958) );
  INV_X2 U5909 ( .A(n5023), .ZN(n5024) );
  INV_X2 U2197 ( .A(n16), .ZN(n814) );
  INV_X2 U1112 ( .A(n1880), .ZN(n813) );
  INV_X2 U4814 ( .A(n4384), .ZN(n4385) );
  AND2_X2 U2426 ( .A1(n2315), .A2(n2314), .ZN(n957) );
  INV_X2 U2158 ( .A(n3975), .ZN(n791) );
  NAND2_X2 U2099 ( .A1(n956), .A2(n3700), .ZN(n4621) );
  INV_X2 U1476 ( .A(n1537), .ZN(n1536) );
  INV_X2 U1598 ( .A(n3088), .ZN(n478) );
  INV_X2 U939 ( .A(n2719), .ZN(n755) );
  INV_X2 U1254 ( .A(n4447), .ZN(n316) );
  INV_X2 U2802 ( .A(n1856), .ZN(n1853) );
  NOR2_X2 U1341 ( .A1(n3057), .A2(n4047), .ZN(n4457) );
  INV_X2 U531 ( .A(n4458), .ZN(n4461) );
  INV_X2 U4809 ( .A(n6674), .ZN(n5227) );
  INV_X2 U1134 ( .A(n2334), .ZN(n261) );
  INV_X2 U1256 ( .A(n2590), .ZN(n5017) );
  INV_X2 U2295 ( .A(n3530), .ZN(n3112) );
  INV_X2 U2991 ( .A(n4870), .ZN(n2627) );
  INV_X2 U1340 ( .A(n4457), .ZN(n348) );
  BUF_X2 U589 ( .A(n4232), .Z(n102) );
  NOR2_X1 U6162 ( .A1(n6027), .A2(n6026), .ZN(n6031) );
  NAND2_X2 U3716 ( .A1(n3889), .A2(n3890), .ZN(n2322) );
  XNOR2_X1 U6146 ( .A(n6026), .B(n6027), .ZN(n5962) );
  INV_X2 U898 ( .A(n3929), .ZN(n1039) );
  INV_X2 U1143 ( .A(n4904), .ZN(n355) );
  INV_X2 U2073 ( .A(n4575), .ZN(n738) );
  INV_X2 U2500 ( .A(n4523), .ZN(n3501) );
  INV_X2 U1731 ( .A(n102), .ZN(n552) );
  NAND2_X2 U3066 ( .A1(n4230), .A2(n1123), .ZN(n4243) );
  NAND2_X2 U1839 ( .A1(n3038), .A2(n3037), .ZN(n2186) );
  NOR2_X2 U1843 ( .A1(n3560), .A2(n4878), .ZN(n3688) );
  INV_X2 U1218 ( .A(n2333), .ZN(n295) );
  INV_X2 U1397 ( .A(n1406), .ZN(n392) );
  INV_X2 U1800 ( .A(n4044), .ZN(n3967) );
  INV_X2 U2742 ( .A(n3985), .ZN(n1173) );
  XNOR2_X1 U6166 ( .A(n6122), .B(n6121), .ZN(n6051) );
  INV_X4 U389 ( .A(n4585), .ZN(n2947) );
  INV_X2 U4706 ( .A(n6201), .ZN(n4262) );
  INV_X1 U2765 ( .A(n4197), .ZN(n4198) );
  INV_X2 U4066 ( .A(n2011), .ZN(n3926) );
  INV_X2 U866 ( .A(n181), .ZN(n273) );
  INV_X2 U1007 ( .A(n3024), .ZN(n447) );
  INV_X2 U2329 ( .A(n1122), .ZN(n905) );
  NAND2_X2 U3375 ( .A1(n1900), .A2(n1901), .ZN(n4255) );
  AOI21_X1 U289 ( .B1(n6114), .B2(n6051), .A(n6112), .ZN(n6054) );
  INV_X2 U213 ( .A(n3898), .ZN(n1498) );
  INV_X2 U1961 ( .A(n3936), .ZN(n768) );
  INV_X2 U223 ( .A(n539), .ZN(n13) );
  NAND2_X2 U4059 ( .A1(n2531), .A2(n3946), .ZN(n4009) );
  NAND2_X2 U1536 ( .A1(n487), .A2(n2598), .ZN(n2599) );
  INV_X2 U972 ( .A(n5210), .ZN(n508) );
  INV_X2 U5585 ( .A(n5685), .ZN(n5686) );
  INV_X2 U1658 ( .A(n1506), .ZN(n507) );
  INV_X2 U825 ( .A(n172), .ZN(n804) );
  NAND2_X2 U2222 ( .A1(n1747), .A2(n3403), .ZN(n834) );
  INV_X2 U2556 ( .A(n3135), .ZN(n5774) );
  INV_X2 U2408 ( .A(n5583), .ZN(n5569) );
  INV_X2 U2690 ( .A(n5691), .ZN(n5684) );
  INV_X2 U2552 ( .A(n5767), .ZN(n1002) );
  INV_X2 U4709 ( .A(n4986), .ZN(n5840) );
  INV_X2 U6089 ( .A(n143), .ZN(n5730) );
  INV_X2 U1227 ( .A(n6423), .ZN(n5740) );
  NAND2_X2 U1863 ( .A1(n2650), .A2(n6348), .ZN(n5813) );
  AND2_X2 U4880 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  NOR2_X2 U2341 ( .A1(n6194), .A2(n5632), .ZN(n5641) );
  INV_X2 U2903 ( .A(b[23]), .ZN(n2569) );
  NAND2_X2 U1246 ( .A1(a[16]), .A2(a[15]), .ZN(n3909) );
  INV_X4 U2640 ( .A(b[12]), .ZN(n3572) );
  XOR2_X2 U2367 ( .A(a[5]), .B(b[12]), .Z(n2706) );
  INV_X4 U109 ( .A(b[0]), .ZN(n4559) );
  INV_X4 U110 ( .A(a[11]), .ZN(n3728) );
  INV_X2 U2881 ( .A(n4784), .ZN(n3203) );
  INV_X2 U2607 ( .A(n4744), .ZN(n1232) );
  NAND2_X2 U5327 ( .A1(a[19]), .A2(n3562), .ZN(n5235) );
  NAND2_X2 U1387 ( .A1(n383), .A2(n384), .ZN(n5365) );
  NAND2_X2 U2399 ( .A1(n3145), .A2(n3144), .ZN(n5231) );
  INV_X2 U2193 ( .A(n5023), .ZN(n810) );
  NOR2_X2 U2144 ( .A1(n2247), .A2(n2250), .ZN(n2246) );
  NOR2_X2 U5069 ( .A1(n4771), .A2(n3324), .ZN(n4802) );
  OR2_X2 U2505 ( .A1(n3055), .A2(n3053), .ZN(n3057) );
  INV_X2 U2129 ( .A(n3616), .ZN(n772) );
  INV_X2 U3618 ( .A(n1489), .ZN(n1488) );
  NAND2_X2 U2593 ( .A1(n3310), .A2(n3309), .ZN(n5237) );
  INV_X2 U2996 ( .A(n3380), .ZN(n2474) );
  INV_X2 U999 ( .A(n3730), .ZN(n1053) );
  INV_X2 U2130 ( .A(n2159), .ZN(n776) );
  OR2_X2 U2501 ( .A1(n5517), .A2(n5516), .ZN(n1679) );
  INV_X2 U2050 ( .A(n41), .ZN(n722) );
  NAND2_X2 U1249 ( .A1(n1488), .A2(n2287), .ZN(n1487) );
  INV_X2 U1643 ( .A(n5451), .ZN(n497) );
  NOR2_X2 U1973 ( .A1(n3277), .A2(n3281), .ZN(n1785) );
  INV_X2 U1897 ( .A(n1482), .ZN(n632) );
  INV_X2 U798 ( .A(n5242), .ZN(n747) );
  INV_X2 U5737 ( .A(n4180), .ZN(n4183) );
  NAND2_X1 U3915 ( .A1(n2355), .A2(n2356), .ZN(n1804) );
  NAND2_X2 U57 ( .A1(n1487), .A2(n3851), .ZN(n3893) );
  INV_X2 U177 ( .A(n3420), .ZN(n3421) );
  INV_X2 U5197 ( .A(n1499), .ZN(n3116) );
  NAND2_X2 U2185 ( .A1(n1925), .A2(n1924), .ZN(n4585) );
  INV_X2 U2083 ( .A(n2813), .ZN(n744) );
  INV_X4 U2736 ( .A(n5421), .ZN(n5434) );
  NOR2_X2 U1864 ( .A1(n4198), .A2(n6378), .ZN(n4201) );
  INV_X2 U2938 ( .A(n4254), .ZN(n1901) );
  XNOR2_X2 U4651 ( .A(n6112), .B(n6117), .ZN(n5964) );
  INV_X2 U336 ( .A(n2576), .ZN(n2881) );
  INV_X4 U2558 ( .A(n1309), .ZN(n5683) );
  INV_X2 U469 ( .A(n5733), .ZN(n64) );
  NOR2_X4 U55 ( .A1(n1590), .A2(n1591), .ZN(n1949) );
  INV_X4 U83 ( .A(n1), .ZN(n4028) );
  INV_X4 U536 ( .A(n2092), .ZN(n88) );
  NAND2_X2 U1784 ( .A1(n1242), .A2(n3313), .ZN(n594) );
  NOR2_X4 U1836 ( .A1(n2950), .A2(n3870), .ZN(n4546) );
  INV_X4 U2909 ( .A(b[19]), .ZN(n3438) );
  INV_X4 U2523 ( .A(b[8]), .ZN(n3342) );
  NOR2_X2 U2247 ( .A1(a[21]), .A2(a[20]), .ZN(n1622) );
  INV_X4 U3373 ( .A(n2889), .ZN(n1326) );
  INV_X4 U95 ( .A(b[2]), .ZN(n2249) );
  NAND3_X2 U145 ( .A1(a[1]), .A2(a[3]), .A3(n4674), .ZN(n4835) );
  NAND2_X2 U1586 ( .A1(n4601), .A2(b[17]), .ZN(n3132) );
  NAND2_X2 U5232 ( .A1(n3507), .A2(a[17]), .ZN(n4767) );
  NOR2_X2 U4505 ( .A1(n2537), .A2(n3540), .ZN(n4029) );
  NOR2_X2 U4667 ( .A1(n465), .A2(n2380), .ZN(n5181) );
  NAND2_X2 U3073 ( .A1(n3052), .A2(n4210), .ZN(n3320) );
  INV_X4 U3981 ( .A(n6459), .ZN(n5079) );
  NAND2_X2 U558 ( .A1(n2794), .A2(n2795), .ZN(n2792) );
  NAND2_X2 U1610 ( .A1(n1740), .A2(n3781), .ZN(n3890) );
  NAND2_X2 U3194 ( .A1(n2103), .A2(n4847), .ZN(n1727) );
  NOR3_X2 U1698 ( .A1(n1736), .A2(n1735), .A3(n1734), .ZN(n3894) );
  NAND2_X2 U3067 ( .A1(n4183), .A2(n4182), .ZN(n4230) );
  NAND2_X2 U1 ( .A1(n2175), .A2(n2174), .ZN(n1975) );
  NOR2_X2 U6 ( .A1(n4123), .A2(n4122), .ZN(n4139) );
  NOR2_X2 U11 ( .A1(n4504), .A2(n2249), .ZN(n3668) );
  NOR3_X2 U22 ( .A1(a[4]), .A2(a[3]), .A3(b[22]), .ZN(n4740) );
  NAND2_X2 U29 ( .A1(n6342), .A2(n6343), .ZN(n2700) );
  INV_X4 U45 ( .A(b[9]), .ZN(n6221) );
  NAND2_X2 U48 ( .A1(a[3]), .A2(b[22]), .ZN(n4700) );
  INV_X4 U59 ( .A(b[22]), .ZN(n566) );
  INV_X8 U65 ( .A(n5895), .ZN(n4829) );
  XNOR2_X2 U84 ( .A(n5720), .B(n5719), .ZN(\d[14]_BAR ) );
  INV_X2 U85 ( .A(n2988), .ZN(n5796) );
  OAI22_X1 U92 ( .A1(n4309), .A2(n4307), .B1(n4305), .B2(n4306), .ZN(n4311) );
  INV_X4 U105 ( .A(n70), .ZN(n396) );
  XNOR2_X1 U107 ( .A(n5832), .B(n5790), .ZN(\d[21]_BAR ) );
  XNOR2_X2 U111 ( .A(n5833), .B(n6164), .ZN(\d[24]_BAR ) );
  NAND2_X1 U115 ( .A1(n806), .A2(b[9]), .ZN(n1456) );
  NOR2_X1 U117 ( .A1(n806), .A2(n2249), .ZN(n2997) );
  NOR2_X1 U121 ( .A1(n806), .A2(n3438), .ZN(n6171) );
  NAND2_X1 U122 ( .A1(n2293), .A2(n3534), .ZN(n2292) );
  INV_X2 U123 ( .A(n2901), .ZN(n6198) );
  INV_X4 U149 ( .A(n6405), .ZN(n529) );
  NAND2_X1 U150 ( .A1(n4844), .A2(n2098), .ZN(n2631) );
  NOR2_X1 U162 ( .A1(b[10]), .A2(n998), .ZN(n2122) );
  INV_X4 U163 ( .A(n2574), .ZN(n3371) );
  INV_X2 U194 ( .A(n2976), .ZN(n3354) );
  INV_X2 U198 ( .A(n5128), .ZN(n5126) );
  INV_X4 U199 ( .A(n6337), .ZN(n5693) );
  INV_X2 U202 ( .A(n1136), .ZN(n179) );
  NOR2_X2 U208 ( .A1(n6339), .A2(n6338), .ZN(n6337) );
  INV_X2 U211 ( .A(n3459), .ZN(n6338) );
  INV_X2 U216 ( .A(n4253), .ZN(n1900) );
  INV_X2 U239 ( .A(n5346), .ZN(n5347) );
  BUF_X4 U249 ( .A(n4160), .Z(n6239) );
  NAND2_X2 U252 ( .A1(n4774), .A2(b[9]), .ZN(n4410) );
  INV_X2 U253 ( .A(n4362), .ZN(n6253) );
  INV_X2 U270 ( .A(n5977), .ZN(n5983) );
  XNOR2_X2 U271 ( .A(n1067), .B(n630), .ZN(n4712) );
  INV_X1 U273 ( .A(n6522), .ZN(n5749) );
  OR2_X4 U275 ( .A1(n2650), .A2(n6348), .ZN(n6453) );
  AND2_X2 U282 ( .A1(n2292), .A2(n2294), .ZN(n6454) );
  INV_X2 U283 ( .A(n1947), .ZN(n6229) );
  NAND2_X2 U286 ( .A1(n5683), .A2(n325), .ZN(n5691) );
  INV_X4 U290 ( .A(n5322), .ZN(n5321) );
  INV_X4 U306 ( .A(n1592), .ZN(n6149) );
  INV_X2 U307 ( .A(n3937), .ZN(n141) );
  NAND2_X2 U314 ( .A1(n1899), .A2(n2553), .ZN(n2552) );
  INV_X2 U317 ( .A(n1416), .ZN(n1415) );
  INV_X2 U338 ( .A(n3707), .ZN(n3706) );
  NAND2_X2 U350 ( .A1(n1007), .A2(n3231), .ZN(n1408) );
  INV_X2 U372 ( .A(n1711), .ZN(n6207) );
  INV_X2 U374 ( .A(n2564), .ZN(n6333) );
  NAND2_X2 U375 ( .A1(n1965), .A2(n1968), .ZN(n2011) );
  NAND2_X2 U376 ( .A1(n128), .A2(n127), .ZN(n1269) );
  NAND2_X2 U377 ( .A1(n6371), .A2(n6372), .ZN(n6374) );
  NAND2_X2 U392 ( .A1(n634), .A2(n633), .ZN(n6351) );
  INV_X2 U403 ( .A(n5289), .ZN(n6150) );
  NAND2_X2 U412 ( .A1(n631), .A2(n632), .ZN(n634) );
  INV_X4 U419 ( .A(n3546), .ZN(n6151) );
  INV_X2 U420 ( .A(n5288), .ZN(n6152) );
  INV_X2 U424 ( .A(n1632), .ZN(n6361) );
  INV_X2 U426 ( .A(n5225), .ZN(n6368) );
  OR2_X2 U427 ( .A1(n1960), .A2(n1255), .ZN(n1254) );
  INV_X2 U431 ( .A(n6316), .ZN(n6448) );
  INV_X2 U435 ( .A(n5064), .ZN(n6153) );
  INV_X2 U439 ( .A(n4455), .ZN(n6237) );
  NOR2_X2 U452 ( .A1(n4341), .A2(n1564), .ZN(n4447) );
  NOR2_X2 U455 ( .A1(n1839), .A2(n1838), .ZN(n4455) );
  INV_X4 U459 ( .A(n6239), .ZN(n4084) );
  BUF_X2 U464 ( .A(n4567), .Z(n6293) );
  INV_X2 U470 ( .A(n2026), .ZN(n6390) );
  INV_X2 U474 ( .A(n4235), .ZN(n3493) );
  XOR2_X2 U496 ( .A(b[8]), .B(a[13]), .Z(n4366) );
  XOR2_X2 U497 ( .A(a[5]), .B(b[9]), .Z(n3796) );
  NAND2_X2 U498 ( .A1(a[23]), .A2(b[22]), .ZN(n6101) );
  XOR2_X2 U503 ( .A(b[7]), .B(a[13]), .Z(n2724) );
  XOR2_X2 U514 ( .A(a[9]), .B(b[3]), .Z(n3993) );
  NOR2_X2 U522 ( .A1(a[5]), .A2(a[6]), .ZN(n6181) );
  XOR2_X2 U542 ( .A(a[3]), .B(b[12]), .Z(n3782) );
  AND2_X2 U543 ( .A1(n3217), .A2(a[9]), .ZN(n962) );
  OR2_X1 U561 ( .A1(n513), .A2(b[18]), .ZN(n6159) );
  NAND2_X1 U566 ( .A1(n4767), .A2(n5293), .ZN(n1195) );
  OAI22_X1 U567 ( .A1(n47), .A2(n3154), .B1(b[23]), .B2(n4797), .ZN(n4799) );
  NAND3_X1 U598 ( .A1(n2569), .A2(a[11]), .A3(n360), .ZN(n5102) );
  NOR2_X1 U599 ( .A1(b[14]), .A2(n5109), .ZN(n4757) );
  INV_X1 U605 ( .A(n6184), .ZN(n3875) );
  NOR2_X1 U613 ( .A1(n4706), .A2(n2889), .ZN(n1792) );
  INV_X2 U616 ( .A(n1445), .ZN(n1439) );
  NOR2_X1 U617 ( .A1(n3300), .A2(n1784), .ZN(n3299) );
  NAND2_X1 U621 ( .A1(n5074), .A2(n4598), .ZN(n2197) );
  INV_X2 U627 ( .A(n4020), .ZN(n350) );
  INV_X2 U633 ( .A(n1483), .ZN(n631) );
  NOR2_X1 U634 ( .A1(n6172), .A2(n6171), .ZN(n6170) );
  NAND3_X1 U639 ( .A1(n2392), .A2(n2439), .A3(n4840), .ZN(n1169) );
  INV_X1 U642 ( .A(n5112), .ZN(n5114) );
  INV_X1 U644 ( .A(n3976), .ZN(n2305) );
  NOR2_X2 U645 ( .A1(n3729), .A2(n4598), .ZN(n159) );
  NOR2_X1 U646 ( .A1(n3780), .A2(n5076), .ZN(n1742) );
  NOR2_X1 U648 ( .A1(n5167), .A2(n5166), .ZN(n1204) );
  INV_X1 U651 ( .A(n5281), .ZN(n2558) );
  NAND2_X1 U653 ( .A1(n5502), .A2(n5503), .ZN(n2068) );
  MUX2_X1 U654 ( .A(n2382), .B(n2510), .S(n566), .Z(n5455) );
  AOI21_X1 U657 ( .B1(n5352), .B2(n5351), .A(n5350), .ZN(n5490) );
  INV_X4 U659 ( .A(b[6]), .ZN(n1324) );
  INV_X1 U666 ( .A(n4628), .ZN(n3340) );
  INV_X2 U668 ( .A(n5252), .ZN(n5256) );
  INV_X2 U669 ( .A(n2539), .ZN(n641) );
  INV_X1 U671 ( .A(n1019), .ZN(n867) );
  NOR2_X1 U672 ( .A1(n6001), .A2(n3164), .ZN(n6003) );
  NAND2_X1 U683 ( .A1(n3211), .A2(n4306), .ZN(n859) );
  NOR2_X1 U684 ( .A1(n5590), .A2(n3164), .ZN(n5587) );
  XNOR2_X1 U694 ( .A(n5778), .B(n5771), .ZN(n5776) );
  INV_X1 U695 ( .A(n3387), .ZN(n3406) );
  NOR2_X1 U706 ( .A1(n5677), .A2(n421), .ZN(n5679) );
  OR2_X1 U717 ( .A1(n465), .A2(n3538), .ZN(n6158) );
  AND2_X4 U718 ( .A1(n758), .A2(b[3]), .ZN(n6160) );
  XOR2_X2 U720 ( .A(a[10]), .B(a[9]), .Z(n6161) );
  INV_X2 U722 ( .A(n4497), .ZN(n189) );
  XOR2_X2 U724 ( .A(a[7]), .B(b[2]), .Z(n6162) );
  INV_X2 U725 ( .A(n4302), .ZN(n1026) );
  XOR2_X2 U727 ( .A(a[11]), .B(b[0]), .Z(n6163) );
  INV_X1 U728 ( .A(n2978), .ZN(n3412) );
  XOR2_X1 U738 ( .A(n1359), .B(n5834), .Z(n6164) );
  XNOR2_X2 U763 ( .A(n4191), .B(n1764), .ZN(n1632) );
  INV_X4 U765 ( .A(n4205), .ZN(n545) );
  NAND2_X2 U766 ( .A1(n1632), .A2(n1116), .ZN(n6363) );
  AOI21_X2 U768 ( .B1(n4205), .B2(n1105), .A(n6178), .ZN(n1770) );
  OAI22_X2 U772 ( .A1(n5221), .A2(n4823), .B1(n4822), .B2(b[23]), .ZN(n4824)
         );
  NOR2_X4 U776 ( .A1(n1121), .A2(a[5]), .ZN(n4823) );
  AOI22_X2 U778 ( .A1(n2412), .A2(n2413), .B1(n1287), .B2(n4321), .ZN(n4323)
         );
  NOR2_X2 U788 ( .A1(n6297), .A2(n2000), .ZN(n2868) );
  INV_X2 U815 ( .A(n3332), .ZN(n6169) );
  NAND2_X2 U820 ( .A1(n2838), .A2(n3939), .ZN(n3626) );
  NAND2_X2 U821 ( .A1(n2011), .A2(n2012), .ZN(n2838) );
  NAND2_X2 U824 ( .A1(n5135), .A2(n6170), .ZN(n1428) );
  NOR2_X2 U830 ( .A1(n2656), .A2(b[19]), .ZN(n6172) );
  NAND2_X2 U858 ( .A1(n6173), .A2(n19), .ZN(n1973) );
  INV_X2 U869 ( .A(n2869), .ZN(n6173) );
  AOI21_X2 U877 ( .B1(n1983), .B2(n1981), .A(n1980), .ZN(n2869) );
  NAND3_X2 U885 ( .A1(n6345), .A2(n4318), .A3(n4319), .ZN(n6174) );
  AOI22_X2 U889 ( .A1(n4601), .A2(b[19]), .B1(n6456), .B2(n3438), .ZN(n1527)
         );
  NAND2_X2 U892 ( .A1(n1415), .A2(n1414), .ZN(n3619) );
  NAND2_X2 U894 ( .A1(n4656), .A2(n4655), .ZN(n3648) );
  AOI21_X2 U895 ( .B1(n3606), .B2(n3605), .A(n4603), .ZN(n4656) );
  AOI22_X2 U906 ( .A1(n2382), .A2(b[11]), .B1(n2510), .B2(n981), .ZN(n1590) );
  NOR2_X2 U908 ( .A1(n1837), .A2(n4290), .ZN(n4301) );
  OAI22_X2 U909 ( .A1(n2286), .A2(n4282), .B1(n2285), .B2(n4281), .ZN(n1837)
         );
  OAI22_X2 U910 ( .A1(n3326), .A2(b[7]), .B1(n3465), .B2(n3581), .ZN(n3237) );
  NOR2_X4 U911 ( .A1(n1000), .A2(n3728), .ZN(n3326) );
  NOR2_X2 U917 ( .A1(n2122), .A2(n6175), .ZN(n2121) );
  INV_X2 U918 ( .A(n6176), .ZN(n6175) );
  NAND2_X2 U924 ( .A1(n440), .A2(b[10]), .ZN(n6176) );
  OAI22_X2 U935 ( .A1(n4050), .A2(n4051), .B1(n6589), .B2(n4049), .ZN(n1839)
         );
  OAI21_X1 U944 ( .B1(n5775), .B2(n3135), .A(n5779), .ZN(n25) );
  NAND2_X2 U945 ( .A1(n2988), .A2(n710), .ZN(n5748) );
  INV_X1 U948 ( .A(n949), .ZN(n6177) );
  INV_X2 U952 ( .A(n6177), .ZN(n6178) );
  AND2_X2 U959 ( .A1(n4171), .A2(n4170), .ZN(n949) );
  INV_X1 U970 ( .A(n6618), .ZN(n4289) );
  INV_X1 U974 ( .A(n2364), .ZN(n6179) );
  INV_X1 U978 ( .A(n6179), .ZN(n6180) );
  NOR2_X4 U979 ( .A1(a[5]), .A2(a[6]), .ZN(n6182) );
  INV_X1 U995 ( .A(n4308), .ZN(n3356) );
  NAND2_X2 U1000 ( .A1(a[1]), .A2(n2563), .ZN(n6183) );
  NAND2_X2 U1001 ( .A1(n4244), .A2(n4243), .ZN(n4307) );
  NAND2_X4 U1012 ( .A1(a[1]), .A2(a[2]), .ZN(n6184) );
  NAND2_X4 U1017 ( .A1(a[1]), .A2(a[2]), .ZN(n6185) );
  INV_X4 U1020 ( .A(n4258), .ZN(n4224) );
  NAND2_X1 U1025 ( .A1(n3405), .A2(n4932), .ZN(n1317) );
  NAND2_X1 U1029 ( .A1(n4886), .A2(n3438), .ZN(n6264) );
  XNOR2_X2 U1035 ( .A(n4102), .B(n1052), .ZN(n1129) );
  NOR3_X4 U1039 ( .A1(n3666), .A2(n3664), .A3(n3665), .ZN(n4102) );
  NAND2_X2 U1043 ( .A1(n2605), .A2(n2606), .ZN(n6186) );
  NAND2_X2 U1058 ( .A1(n1151), .A2(n396), .ZN(n6187) );
  INV_X2 U1059 ( .A(n845), .ZN(n6188) );
  INV_X2 U1061 ( .A(n4635), .ZN(n2905) );
  XNOR2_X2 U1062 ( .A(n5820), .B(n6189), .ZN(\d[23]_BAR ) );
  NAND2_X1 U1080 ( .A1(n1324), .A2(n1060), .ZN(n3741) );
  OAI21_X1 U1087 ( .B1(n2792), .B2(n4564), .A(n4612), .ZN(n2013) );
  NAND2_X2 U1096 ( .A1(n4032), .A2(n4031), .ZN(n6191) );
  XNOR2_X2 U1113 ( .A(n5826), .B(n5825), .ZN(\d[22]_BAR ) );
  NAND2_X2 U1151 ( .A1(n872), .A2(n871), .ZN(n5260) );
  INV_X2 U1152 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U1163 ( .A1(n1013), .A2(n1902), .ZN(n6194) );
  NOR2_X2 U1180 ( .A1(n4716), .A2(n4712), .ZN(n1144) );
  AND2_X2 U1189 ( .A1(n3506), .A2(n4422), .ZN(n309) );
  NAND2_X1 U1194 ( .A1(n5454), .A2(b[22]), .ZN(n223) );
  INV_X8 U1195 ( .A(a[3]), .ZN(n4492) );
  INV_X8 U1197 ( .A(a[3]), .ZN(n1066) );
  INV_X2 U1205 ( .A(n3073), .ZN(n2692) );
  INV_X1 U1211 ( .A(n4654), .ZN(n1069) );
  NAND3_X1 U1220 ( .A1(n4079), .A2(n4009), .A3(n1257), .ZN(n3589) );
  NAND2_X1 U1228 ( .A1(n5373), .A2(n2977), .ZN(n927) );
  NAND2_X2 U1251 ( .A1(n2310), .A2(n1298), .ZN(n1294) );
  INV_X2 U1263 ( .A(n2544), .ZN(n836) );
  INV_X2 U1282 ( .A(n5069), .ZN(n1378) );
  NAND2_X2 U1307 ( .A1(n6184), .A2(a[3]), .ZN(n3772) );
  NAND2_X2 U1308 ( .A1(n1266), .A2(n1264), .ZN(n6199) );
  NAND2_X2 U1311 ( .A1(n1266), .A2(n1264), .ZN(n3596) );
  INV_X2 U1313 ( .A(n1771), .ZN(n6371) );
  NAND3_X2 U1314 ( .A1(n340), .A2(n2218), .A3(n4918), .ZN(n6200) );
  XNOR2_X1 U1316 ( .A(n1126), .B(n4227), .ZN(n6201) );
  NAND2_X1 U1333 ( .A1(n1181), .A2(n1182), .ZN(n6202) );
  NOR2_X4 U1336 ( .A1(n4224), .A2(n4256), .ZN(n1126) );
  NAND3_X2 U1337 ( .A1(n3826), .A2(a[10]), .A3(a[9]), .ZN(n4887) );
  NOR2_X1 U1343 ( .A1(n5895), .A2(n3572), .ZN(n3300) );
  NAND2_X1 U1344 ( .A1(n5895), .A2(b[1]), .ZN(n1645) );
  NAND3_X2 U1347 ( .A1(a[6]), .A2(a[5]), .A3(n4689), .ZN(n6203) );
  NAND2_X4 U1349 ( .A1(n1443), .A2(n1444), .ZN(n4883) );
  OAI21_X1 U1353 ( .B1(n4981), .B2(n5094), .A(n343), .ZN(n6205) );
  OAI21_X1 U1354 ( .B1(n4981), .B2(n5094), .A(n343), .ZN(n5380) );
  NAND3_X2 U1356 ( .A1(n1690), .A2(n1840), .A3(n2266), .ZN(n6206) );
  INV_X2 U1358 ( .A(n2030), .ZN(n1447) );
  INV_X1 U1377 ( .A(n1711), .ZN(n4869) );
  NAND2_X1 U1400 ( .A1(n1786), .A2(n4867), .ZN(n6209) );
  INV_X2 U1408 ( .A(n1591), .ZN(n1588) );
  NAND2_X1 U1412 ( .A1(n5162), .A2(n2422), .ZN(n6210) );
  NOR2_X1 U1420 ( .A1(a[3]), .A2(n365), .ZN(n6212) );
  NOR2_X1 U1441 ( .A1(b[12]), .A2(n5473), .ZN(n1784) );
  NOR2_X4 U1454 ( .A1(n1064), .A2(n1066), .ZN(n2129) );
  OAI21_X1 U1457 ( .B1(n4029), .B2(n4028), .A(n3618), .ZN(n6216) );
  AOI21_X2 U1460 ( .B1(n4879), .B2(n2827), .A(n3687), .ZN(n3686) );
  NAND2_X2 U1463 ( .A1(n6220), .A2(n6219), .ZN(n3787) );
  NAND2_X1 U1464 ( .A1(b[9]), .A2(n4601), .ZN(n6219) );
  NAND2_X2 U1470 ( .A1(n3614), .A2(n6221), .ZN(n6220) );
  NAND3_X2 U1471 ( .A1(n1272), .A2(n1270), .A3(n1273), .ZN(n6222) );
  NAND3_X2 U1473 ( .A1(n6223), .A2(n2417), .A3(n2414), .ZN(n2468) );
  NAND3_X2 U1475 ( .A1(n2416), .A2(n1807), .A3(n2418), .ZN(n6223) );
  NAND2_X2 U1489 ( .A1(n1624), .A2(n6224), .ZN(n1625) );
  NOR2_X2 U1490 ( .A1(n6226), .A2(n6225), .ZN(n6224) );
  NOR2_X2 U1497 ( .A1(n2513), .A2(n5007), .ZN(n6225) );
  NOR2_X2 U1500 ( .A1(n1895), .A2(n5006), .ZN(n6226) );
  NAND3_X2 U1505 ( .A1(n2608), .A2(n4579), .A3(n2612), .ZN(n6291) );
  NAND3_X2 U1526 ( .A1(n2154), .A2(n5325), .A3(n6092), .ZN(n2153) );
  NOR2_X2 U1527 ( .A1(n5834), .A2(n2087), .ZN(n5325) );
  INV_X4 U1528 ( .A(n3106), .ZN(n514) );
  OAI22_X2 U1529 ( .A1(n6228), .A2(n1048), .B1(n5285), .B2(n5284), .ZN(n5355)
         );
  NOR2_X2 U1530 ( .A1(n5282), .A2(n1037), .ZN(n6228) );
  NAND2_X2 U1541 ( .A1(n226), .A2(n225), .ZN(n3319) );
  NAND2_X2 U1543 ( .A1(n3273), .A2(n1485), .ZN(n225) );
  NAND2_X2 U1544 ( .A1(n3628), .A2(n3107), .ZN(n6256) );
  NAND2_X2 U1545 ( .A1(n514), .A2(n3627), .ZN(n3628) );
  NOR2_X2 U1556 ( .A1(n6229), .A2(n6422), .ZN(n3477) );
  NAND2_X2 U1565 ( .A1(n6230), .A2(n4934), .ZN(n1750) );
  INV_X2 U1566 ( .A(n4931), .ZN(n6230) );
  AOI22_X2 U1573 ( .A1(n6231), .A2(n6159), .B1(n2702), .B2(n4933), .ZN(n1215)
         );
  AOI22_X2 U1592 ( .A1(n4610), .A2(b[7]), .B1(n3465), .B2(n4609), .ZN(n3868)
         );
  NAND2_X4 U1605 ( .A1(n6188), .A2(n3058), .ZN(n4610) );
  NAND2_X2 U1622 ( .A1(n2294), .A2(n2237), .ZN(n2236) );
  NAND2_X2 U1638 ( .A1(n6232), .A2(n270), .ZN(n4300) );
  NAND2_X2 U1639 ( .A1(n268), .A2(n269), .ZN(n6232) );
  INV_X4 U1641 ( .A(n4294), .ZN(n4005) );
  NAND2_X2 U1642 ( .A1(n3989), .A2(n6233), .ZN(n3998) );
  NOR2_X2 U1662 ( .A1(n6235), .A2(n6234), .ZN(n6233) );
  NOR2_X2 U1667 ( .A1(n4217), .A2(b[10]), .ZN(n6235) );
  NAND2_X2 U1669 ( .A1(n3746), .A2(n3948), .ZN(n3120) );
  NAND2_X2 U1670 ( .A1(n6236), .A2(n542), .ZN(n2093) );
  NAND2_X2 U1678 ( .A1(n540), .A2(n541), .ZN(n6236) );
  NOR2_X2 U1696 ( .A1(n6157), .A2(n4173), .ZN(n1116) );
  OAI22_X2 U1713 ( .A1(n1847), .A2(b[22]), .B1(n2244), .B2(n5105), .ZN(n2056)
         );
  NAND3_X4 U1715 ( .A1(n2162), .A2(a[5]), .A3(a[6]), .ZN(n2244) );
  NAND2_X2 U1716 ( .A1(n6237), .A2(n4456), .ZN(n1776) );
  NAND2_X2 U1720 ( .A1(n1839), .A2(n1838), .ZN(n4456) );
  NAND2_X2 U1721 ( .A1(n6238), .A2(n546), .ZN(n4203) );
  NAND2_X2 U1723 ( .A1(n544), .A2(n545), .ZN(n6238) );
  NOR2_X2 U1732 ( .A1(n6240), .A2(n2873), .ZN(n2871) );
  INV_X2 U1742 ( .A(n5340), .ZN(n6240) );
  NOR2_X2 U1743 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  NOR2_X1 U1749 ( .A1(n5076), .A2(b[4]), .ZN(n4054) );
  NAND2_X2 U1756 ( .A1(n6241), .A2(n499), .ZN(n5348) );
  NAND2_X2 U1758 ( .A1(n498), .A2(n497), .ZN(n6241) );
  NOR2_X2 U1760 ( .A1(n6245), .A2(n6243), .ZN(n6242) );
  NOR2_X2 U1780 ( .A1(n3431), .A2(b[4]), .ZN(n6245) );
  NAND2_X2 U1782 ( .A1(n6246), .A2(n769), .ZN(n2189) );
  NAND2_X2 U1786 ( .A1(n767), .A2(n768), .ZN(n6246) );
  NAND3_X1 U1792 ( .A1(n5380), .A2(n2278), .A3(n2782), .ZN(n2781) );
  NAND2_X2 U1824 ( .A1(n6249), .A2(n426), .ZN(n429) );
  INV_X2 U1827 ( .A(n1541), .ZN(n6249) );
  NOR2_X2 U1831 ( .A1(n1536), .A2(n425), .ZN(n1541) );
  NAND2_X2 U1832 ( .A1(n6250), .A2(n2444), .ZN(n3930) );
  OAI21_X2 U1840 ( .B1(n2443), .B2(n3621), .A(n3929), .ZN(n6250) );
  AOI21_X2 U1842 ( .B1(n3940), .B2(n2838), .A(n3939), .ZN(n1416) );
  NOR2_X2 U1853 ( .A1(n2778), .A2(n2785), .ZN(n3678) );
  NAND2_X2 U1896 ( .A1(n1056), .A2(n3911), .ZN(n1293) );
  AOI21_X2 U1906 ( .B1(n4931), .B2(n4212), .A(n3540), .ZN(n2602) );
  NAND3_X1 U1907 ( .A1(n2378), .A2(n4045), .A3(n4998), .ZN(n4212) );
  NAND2_X2 U1913 ( .A1(n6252), .A2(n764), .ZN(n1593) );
  NAND2_X2 U1914 ( .A1(n762), .A2(n763), .ZN(n6252) );
  INV_X4 U1918 ( .A(n6437), .ZN(n6436) );
  NAND2_X2 U1921 ( .A1(n6253), .A2(n4014), .ZN(n2926) );
  NAND2_X4 U1925 ( .A1(a[11]), .A2(a[12]), .ZN(n4362) );
  NAND2_X2 U1926 ( .A1(n6254), .A2(n6403), .ZN(n5085) );
  NAND2_X2 U1929 ( .A1(n125), .A2(n5084), .ZN(n6254) );
  NAND2_X2 U1934 ( .A1(n6255), .A2(n6385), .ZN(n2651) );
  NAND3_X2 U1958 ( .A1(n1047), .A2(n3095), .A3(n120), .ZN(n6255) );
  NAND2_X2 U1959 ( .A1(n6256), .A2(n3629), .ZN(n3525) );
  INV_X4 U1962 ( .A(n2327), .ZN(n2326) );
  NAND2_X4 U1965 ( .A1(n361), .A2(n468), .ZN(n2327) );
  INV_X2 U1976 ( .A(n4380), .ZN(n2991) );
  NAND2_X2 U1978 ( .A1(n4020), .A2(n4019), .ZN(n4380) );
  AOI22_X2 U1983 ( .A1(n6258), .A2(n4803), .B1(n4802), .B2(n400), .ZN(n4804)
         );
  NAND2_X2 U1998 ( .A1(n6260), .A2(n6259), .ZN(n6258) );
  NAND2_X2 U2007 ( .A1(n1837), .A2(n4290), .ZN(n1836) );
  NAND2_X4 U2008 ( .A1(n3405), .A2(n3829), .ZN(n3832) );
  NOR2_X4 U2020 ( .A1(n1201), .A2(n4301), .ZN(n4303) );
  NAND2_X2 U2023 ( .A1(n2313), .A2(n2978), .ZN(n2312) );
  NAND3_X2 U2024 ( .A1(n2526), .A2(n2525), .A3(n2527), .ZN(n2978) );
  AOI22_X2 U2026 ( .A1(n6221), .A2(n3230), .B1(n5136), .B2(b[9]), .ZN(n3575)
         );
  AOI21_X2 U2040 ( .B1(n5177), .B2(n5176), .A(n3384), .ZN(n5259) );
  INV_X4 U2059 ( .A(n5206), .ZN(n3499) );
  INV_X2 U2086 ( .A(n5113), .ZN(n3449) );
  BUF_X4 U2116 ( .A(n1888), .Z(n6263) );
  AOI22_X2 U2118 ( .A1(n6265), .A2(n6264), .B1(n2701), .B2(n2326), .ZN(n4920)
         );
  NAND2_X2 U2119 ( .A1(n6439), .A2(b[19]), .ZN(n6265) );
  AOI22_X2 U2120 ( .A1(n6266), .A2(n3030), .B1(n3029), .B2(n3832), .ZN(n3843)
         );
  NOR2_X2 U2123 ( .A1(n439), .A2(n3033), .ZN(n6266) );
  OAI22_X2 U2124 ( .A1(n2619), .A2(n2615), .B1(n2614), .B2(n6267), .ZN(n4519)
         );
  NAND2_X2 U2127 ( .A1(n4517), .A2(n4518), .ZN(n6267) );
  NAND2_X2 U2133 ( .A1(n5156), .A2(n5157), .ZN(n5158) );
  NAND2_X2 U2140 ( .A1(n1541), .A2(n4108), .ZN(n428) );
  XNOR2_X2 U2149 ( .A(n4624), .B(n4622), .ZN(n1366) );
  NAND2_X2 U2152 ( .A1(n3084), .A2(n2372), .ZN(n4622) );
  NAND2_X1 U2169 ( .A1(n558), .A2(b[11]), .ZN(n6450) );
  INV_X4 U2174 ( .A(n6268), .ZN(n122) );
  NOR2_X2 U2176 ( .A1(n2173), .A2(n4300), .ZN(n6268) );
  NAND2_X2 U2189 ( .A1(n6269), .A2(n4891), .ZN(n1660) );
  NAND2_X2 U2190 ( .A1(n495), .A2(n494), .ZN(n6269) );
  NAND2_X2 U2194 ( .A1(n6270), .A2(n293), .ZN(n2082) );
  NAND2_X2 U2215 ( .A1(n4178), .A2(n6272), .ZN(n4181) );
  NOR2_X2 U2218 ( .A1(n6274), .A2(n6273), .ZN(n6272) );
  NOR2_X2 U2219 ( .A1(n4216), .A2(n3465), .ZN(n6273) );
  NOR2_X2 U2226 ( .A1(n4217), .A2(b[7]), .ZN(n6274) );
  OAI21_X1 U2234 ( .B1(n3405), .B2(n2737), .A(n4696), .ZN(n1576) );
  BUF_X4 U2238 ( .A(n2827), .Z(n1499) );
  NAND3_X2 U2240 ( .A1(n4738), .A2(n4739), .A3(n4737), .ZN(n1544) );
  NAND3_X2 U2248 ( .A1(n6276), .A2(n6275), .A3(n2452), .ZN(n6277) );
  INV_X2 U2258 ( .A(n4765), .ZN(n6276) );
  INV_X2 U2259 ( .A(n3078), .ZN(n97) );
  NAND3_X2 U2265 ( .A1(n2174), .A2(n2175), .A3(n1977), .ZN(n3078) );
  NAND2_X2 U2280 ( .A1(n2635), .A2(n1146), .ZN(n2802) );
  NAND2_X2 U2287 ( .A1(n4696), .A2(n2737), .ZN(n1167) );
  NAND3_X2 U2291 ( .A1(n3026), .A2(n633), .A3(n634), .ZN(n4737) );
  NAND2_X2 U2294 ( .A1(n6590), .A2(n4975), .ZN(n3466) );
  NAND2_X2 U2302 ( .A1(n2020), .A2(n6468), .ZN(n4975) );
  NAND2_X2 U2303 ( .A1(n1141), .A2(n6278), .ZN(n4476) );
  OAI21_X1 U2305 ( .B1(n4388), .B2(n4387), .A(n3229), .ZN(n6278) );
  NAND2_X2 U2306 ( .A1(n3156), .A2(n1059), .ZN(n3094) );
  NAND2_X2 U2308 ( .A1(n2021), .A2(n1305), .ZN(n2949) );
  INV_X2 U2315 ( .A(n3414), .ZN(n6279) );
  OR2_X2 U2342 ( .A1(n6015), .A2(n4982), .ZN(n997) );
  NOR2_X2 U2349 ( .A1(n5381), .A2(n6205), .ZN(n6015) );
  NAND2_X2 U2363 ( .A1(n860), .A2(n859), .ZN(n4267) );
  NAND2_X2 U2365 ( .A1(n6283), .A2(n2839), .ZN(n1436) );
  NAND2_X2 U2370 ( .A1(n2841), .A2(n2842), .ZN(n6283) );
  INV_X4 U2377 ( .A(n1465), .ZN(n2765) );
  NAND3_X2 U2416 ( .A1(n2768), .A2(n5976), .A3(n5919), .ZN(n5864) );
  NAND2_X2 U2428 ( .A1(n2215), .A2(n3648), .ZN(n6284) );
  NOR2_X2 U2438 ( .A1(n2623), .A2(n2622), .ZN(n6286) );
  NAND2_X2 U2457 ( .A1(n2929), .A2(n3409), .ZN(n3574) );
  NAND3_X2 U2461 ( .A1(n1381), .A2(n4871), .A3(n1380), .ZN(n2929) );
  NAND2_X2 U2462 ( .A1(n6287), .A2(n2482), .ZN(n2939) );
  NOR2_X2 U2463 ( .A1(n4519), .A2(n4520), .ZN(n4574) );
  NAND2_X2 U2468 ( .A1(n2790), .A2(n2788), .ZN(n4520) );
  NAND2_X2 U2482 ( .A1(n191), .A2(n692), .ZN(n6289) );
  NAND2_X2 U2507 ( .A1(n6290), .A2(n4553), .ZN(n1259) );
  NAND2_X2 U2515 ( .A1(n2938), .A2(n2937), .ZN(n6290) );
  AOI22_X2 U2527 ( .A1(n3591), .A2(n3592), .B1(n3777), .B2(n4408), .ZN(n3802)
         );
  NAND2_X4 U2528 ( .A1(n2609), .A2(n6291), .ZN(n3492) );
  NAND2_X2 U2533 ( .A1(n1272), .A2(n1273), .ZN(n128) );
  NOR2_X2 U2536 ( .A1(n1045), .A2(n5005), .ZN(n1517) );
  NAND2_X2 U2544 ( .A1(n6294), .A2(n352), .ZN(n3973) );
  NAND2_X2 U2545 ( .A1(n350), .A2(n351), .ZN(n6294) );
  NAND2_X1 U2548 ( .A1(n495), .A2(n494), .ZN(n436) );
  NAND2_X2 U2584 ( .A1(n492), .A2(n493), .ZN(n495) );
  INV_X2 U2591 ( .A(n6295), .ZN(n1256) );
  NOR2_X1 U2597 ( .A1(n1215), .A2(n4836), .ZN(n6295) );
  NAND2_X2 U2601 ( .A1(n2190), .A2(n2191), .ZN(n2066) );
  NAND2_X2 U2605 ( .A1(n1184), .A2(n1043), .ZN(n2913) );
  INV_X4 U2608 ( .A(n6296), .ZN(n3634) );
  NAND2_X2 U2611 ( .A1(n3529), .A2(n3528), .ZN(n6296) );
  AOI22_X2 U2622 ( .A1(n2382), .A2(b[5]), .B1(n2510), .B2(n3870), .ZN(n6297)
         );
  NAND3_X2 U2628 ( .A1(n2572), .A2(n2571), .A3(n1795), .ZN(n1518) );
  NAND2_X2 U2631 ( .A1(n1250), .A2(n2888), .ZN(n2572) );
  INV_X4 U2638 ( .A(n6298), .ZN(n4521) );
  NAND2_X2 U2646 ( .A1(n4412), .A2(n4413), .ZN(n6298) );
  AOI21_X2 U2648 ( .B1(n2658), .B2(n4964), .A(n4963), .ZN(n5032) );
  NAND3_X2 U2663 ( .A1(n1480), .A2(n209), .A3(n1478), .ZN(n2658) );
  NAND2_X2 U2672 ( .A1(n6365), .A2(n2911), .ZN(n451) );
  INV_X2 U2678 ( .A(n6299), .ZN(n1357) );
  NAND2_X2 U2681 ( .A1(n628), .A2(n6601), .ZN(n6299) );
  NOR2_X2 U2707 ( .A1(n1915), .A2(n5662), .ZN(n5666) );
  NAND2_X4 U2723 ( .A1(n876), .A2(n875), .ZN(n1915) );
  NAND2_X2 U2724 ( .A1(n5805), .A2(n3672), .ZN(n2381) );
  AOI22_X2 U2759 ( .A1(n3217), .A2(n2656), .B1(n806), .B2(b[17]), .ZN(n5005)
         );
  NAND2_X2 U2776 ( .A1(n1111), .A2(n118), .ZN(n4769) );
  NAND2_X2 U2779 ( .A1(n2303), .A2(n557), .ZN(n5012) );
  NAND2_X2 U2806 ( .A1(n336), .A2(n335), .ZN(n2373) );
  NAND2_X2 U2809 ( .A1(n1682), .A2(n2447), .ZN(n2446) );
  NAND2_X2 U2831 ( .A1(n6569), .A2(n435), .ZN(n4545) );
  INV_X2 U2833 ( .A(n3335), .ZN(n2943) );
  XNOR2_X2 U2848 ( .A(n1366), .B(n1040), .ZN(n3335) );
  NAND2_X2 U2857 ( .A1(n6300), .A2(n287), .ZN(n23) );
  INV_X2 U2858 ( .A(n2550), .ZN(n6300) );
  NAND2_X2 U2860 ( .A1(n1871), .A2(n4247), .ZN(n2550) );
  NAND2_X2 U2891 ( .A1(n6302), .A2(n6301), .ZN(n1525) );
  NAND2_X2 U2898 ( .A1(n6326), .A2(n3465), .ZN(n6301) );
  NAND2_X2 U2900 ( .A1(b[7]), .A2(n760), .ZN(n6302) );
  NOR3_X2 U2914 ( .A1(n1920), .A2(n1921), .A3(n1919), .ZN(n4103) );
  NOR2_X2 U2923 ( .A1(n4874), .A2(n1949), .ZN(n4877) );
  NAND2_X2 U2931 ( .A1(n6303), .A2(n790), .ZN(n2416) );
  NAND2_X2 U2948 ( .A1(n6304), .A2(n4330), .ZN(n4333) );
  NAND2_X2 U2972 ( .A1(n6418), .A2(n2128), .ZN(n4328) );
  NAND2_X2 U2990 ( .A1(n3212), .A2(n6305), .ZN(n3211) );
  NAND3_X2 U2992 ( .A1(n3355), .A2(n4307), .A3(n4308), .ZN(n6305) );
  NAND2_X4 U2993 ( .A1(n6306), .A2(n1276), .ZN(n4612) );
  NAND2_X2 U3000 ( .A1(n87), .A2(n3081), .ZN(n6306) );
  INV_X4 U3001 ( .A(n4453), .ZN(n6404) );
  NAND2_X2 U3004 ( .A1(n4578), .A2(n4577), .ZN(n1712) );
  NAND2_X2 U3008 ( .A1(n119), .A2(n739), .ZN(n4578) );
  NAND2_X2 U3024 ( .A1(n6307), .A2(n863), .ZN(n4305) );
  NAND2_X2 U3030 ( .A1(n861), .A2(n862), .ZN(n6307) );
  NAND2_X2 U3034 ( .A1(n6407), .A2(n6308), .ZN(n3026) );
  NAND4_X1 U3044 ( .A1(n993), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(n6308)
         );
  INV_X2 U3051 ( .A(n6309), .ZN(n2043) );
  NAND2_X2 U3056 ( .A1(n812), .A2(n811), .ZN(n6309) );
  NAND3_X2 U3063 ( .A1(n3903), .A2(n3746), .A3(n3902), .ZN(n3707) );
  NAND2_X2 U3071 ( .A1(n3021), .A2(n3016), .ZN(n2126) );
  NOR3_X2 U3078 ( .A1(n6310), .A2(n3433), .A3(n3432), .ZN(n4550) );
  NOR3_X2 U3092 ( .A1(n3435), .A2(n3436), .A3(n3437), .ZN(n6310) );
  NAND2_X2 U3103 ( .A1(n454), .A2(n6431), .ZN(n6311) );
  NOR2_X2 U3182 ( .A1(n4217), .A2(b[8]), .ZN(n1349) );
  NAND2_X2 U3184 ( .A1(n1039), .A2(n3928), .ZN(n2010) );
  NAND2_X2 U3192 ( .A1(n3495), .A2(n2993), .ZN(n364) );
  AOI22_X2 U3193 ( .A1(n2382), .A2(b[15]), .B1(n2510), .B2(n984), .ZN(n3531)
         );
  NAND2_X2 U3217 ( .A1(n517), .A2(n6315), .ZN(n1658) );
  NAND2_X2 U3221 ( .A1(n3627), .A2(n3106), .ZN(n6315) );
  NAND2_X2 U3230 ( .A1(n4368), .A2(n3067), .ZN(n6316) );
  INV_X4 U3245 ( .A(n6317), .ZN(n5176) );
  NOR2_X2 U3251 ( .A1(n5116), .A2(n5115), .ZN(n6317) );
  NOR2_X2 U3252 ( .A1(n4383), .A2(n4384), .ZN(n3017) );
  NAND2_X2 U3254 ( .A1(n6319), .A2(n6318), .ZN(n3852) );
  NAND2_X2 U3258 ( .A1(n4506), .A2(b[10]), .ZN(n6319) );
  NAND2_X2 U3263 ( .A1(n4728), .A2(n1132), .ZN(n2736) );
  NAND2_X2 U3267 ( .A1(n6320), .A2(n176), .ZN(n2810) );
  INV_X2 U3268 ( .A(n5304), .ZN(n6320) );
  NAND2_X2 U3274 ( .A1(n244), .A2(n746), .ZN(n5304) );
  OAI21_X2 U3290 ( .B1(n5074), .B2(b[16]), .A(n6321), .ZN(n2036) );
  NAND2_X2 U3301 ( .A1(n6322), .A2(b[16]), .ZN(n6321) );
  AOI21_X2 U3317 ( .B1(n1225), .B2(n3778), .A(n1051), .ZN(n1512) );
  NOR2_X2 U3340 ( .A1(n3788), .A2(n414), .ZN(n3789) );
  INV_X1 U3345 ( .A(n1030), .ZN(n3221) );
  AOI22_X1 U3351 ( .A1(n2904), .A2(n2905), .B1(n4635), .B2(n4637), .ZN(n2538)
         );
  NAND2_X4 U3360 ( .A1(n3709), .A2(n6474), .ZN(n3067) );
  NOR3_X4 U3392 ( .A1(n3298), .A2(a[16]), .A3(a[15]), .ZN(n6326) );
  INV_X8 U3402 ( .A(a[17]), .ZN(n3298) );
  NAND2_X2 U3403 ( .A1(n1504), .A2(n192), .ZN(n6327) );
  INV_X4 U3410 ( .A(n193), .ZN(n192) );
  INV_X2 U3416 ( .A(n3554), .ZN(n269) );
  OR2_X2 U3428 ( .A1(n3799), .A2(n4002), .ZN(n965) );
  NOR2_X4 U3438 ( .A1(n3396), .A2(n5729), .ZN(n473) );
  OAI21_X2 U3441 ( .B1(b[21]), .B2(n3586), .A(n3587), .ZN(n5050) );
  NAND2_X1 U3443 ( .A1(n328), .A2(n3538), .ZN(n2618) );
  NAND2_X2 U3446 ( .A1(n2710), .A2(n4933), .ZN(n3533) );
  NOR2_X4 U3447 ( .A1(a[22]), .A2(a[21]), .ZN(n6328) );
  OAI21_X2 U3459 ( .B1(n3134), .B2(n3149), .A(n3220), .ZN(n6329) );
  NAND2_X2 U3473 ( .A1(n133), .A2(n3109), .ZN(n6330) );
  NAND2_X2 U3475 ( .A1(n834), .A2(n835), .ZN(n6331) );
  OAI21_X1 U3480 ( .B1(n2366), .B2(n3347), .A(n4471), .ZN(n2365) );
  NAND2_X1 U3483 ( .A1(n4940), .A2(n6221), .ZN(n4411) );
  NAND2_X1 U3484 ( .A1(n981), .A2(n4940), .ZN(n1457) );
  NAND2_X4 U3491 ( .A1(n591), .A2(n590), .ZN(n4668) );
  NAND2_X2 U3502 ( .A1(n4445), .A2(n3604), .ZN(n579) );
  OAI22_X2 U3506 ( .A1(n4444), .A2(n6448), .B1(n4368), .B2(n3067), .ZN(n4371)
         );
  NAND2_X4 U3526 ( .A1(n1497), .A2(n1494), .ZN(n4314) );
  NAND2_X1 U3527 ( .A1(n4199), .A2(n2564), .ZN(n6334) );
  NAND2_X2 U3537 ( .A1(n775), .A2(n774), .ZN(n4199) );
  INV_X2 U3538 ( .A(n5665), .ZN(n4153) );
  NOR2_X1 U3556 ( .A1(n5136), .A2(n3342), .ZN(n2252) );
  INV_X2 U3558 ( .A(n4504), .ZN(n4337) );
  NOR2_X1 U3583 ( .A1(n1215), .A2(n3294), .ZN(n3503) );
  INV_X2 U3590 ( .A(n2335), .ZN(n4083) );
  NOR2_X4 U3591 ( .A1(n5164), .A2(n5165), .ZN(n2074) );
  NAND2_X2 U3597 ( .A1(n3456), .A2(n3454), .ZN(n6339) );
  NAND2_X1 U3611 ( .A1(n3902), .A2(n266), .ZN(n3948) );
  NAND2_X1 U3624 ( .A1(n4544), .A2(a[23]), .ZN(n4561) );
  INV_X2 U3634 ( .A(n3842), .ZN(n3845) );
  NAND2_X4 U3643 ( .A1(n885), .A2(n886), .ZN(n5258) );
  NAND2_X2 U3644 ( .A1(a[5]), .A2(a[6]), .ZN(n6342) );
  INV_X4 U3656 ( .A(a[5]), .ZN(n6340) );
  INV_X8 U3667 ( .A(a[6]), .ZN(n6341) );
  NOR2_X2 U3668 ( .A1(n3962), .A2(n2700), .ZN(n3904) );
  NAND2_X1 U3688 ( .A1(n3265), .A2(n909), .ZN(n6344) );
  NAND2_X2 U3689 ( .A1(n2160), .A2(n4322), .ZN(n6345) );
  INV_X4 U3690 ( .A(n4323), .ZN(n2160) );
  NAND2_X2 U3692 ( .A1(n5899), .A2(b[11]), .ZN(n134) );
  OAI21_X1 U3694 ( .B1(n5899), .B2(n1884), .A(n1061), .ZN(n1219) );
  INV_X8 U3703 ( .A(n3512), .ZN(n5899) );
  XNOR2_X2 U3712 ( .A(n6346), .B(b[1]), .ZN(n2733) );
  INV_X8 U3717 ( .A(a[19]), .ZN(n6346) );
  INV_X2 U3719 ( .A(n4736), .ZN(n560) );
  INV_X1 U3725 ( .A(n2374), .ZN(n6347) );
  INV_X2 U3742 ( .A(n6347), .ZN(n6348) );
  NAND2_X4 U3743 ( .A1(n4928), .A2(n433), .ZN(n5027) );
  NAND2_X1 U3744 ( .A1(n1107), .A2(n3438), .ZN(n116) );
  NOR2_X2 U3749 ( .A1(n2776), .A2(n5526), .ZN(n4436) );
  OAI21_X1 U3750 ( .B1(n5026), .B2(n5025), .A(n2751), .ZN(n5028) );
  NAND2_X2 U3751 ( .A1(n1948), .A2(n1947), .ZN(n6349) );
  NAND2_X2 U3758 ( .A1(n1948), .A2(n1947), .ZN(n2532) );
  INV_X2 U3765 ( .A(n2538), .ZN(n640) );
  NAND2_X2 U3770 ( .A1(n3477), .A2(n5093), .ZN(n6350) );
  NAND2_X1 U3782 ( .A1(n4893), .A2(n1531), .ZN(n3196) );
  AOI22_X1 U3783 ( .A1(n4705), .A2(b[15]), .B1(n984), .B2(n998), .ZN(n1793) );
  XNOR2_X2 U3797 ( .A(a[15]), .B(b[22]), .ZN(n5220) );
  INV_X8 U3805 ( .A(b[22]), .ZN(n5105) );
  XNOR2_X2 U3816 ( .A(a[1]), .B(b[22]), .ZN(n4418) );
  XNOR2_X2 U3850 ( .A(a[11]), .B(b[22]), .ZN(n4997) );
  INV_X1 U3857 ( .A(n3404), .ZN(n6352) );
  INV_X2 U3864 ( .A(n6352), .ZN(n6353) );
  INV_X1 U3865 ( .A(n1461), .ZN(n5161) );
  INV_X2 U3873 ( .A(n1467), .ZN(n663) );
  NAND2_X2 U3878 ( .A1(n2195), .A2(n3887), .ZN(n1403) );
  NOR2_X4 U3885 ( .A1(n2194), .A2(n3228), .ZN(n2437) );
  NAND2_X1 U3886 ( .A1(n5062), .A2(n5064), .ZN(n6355) );
  NAND2_X2 U3887 ( .A1(n6354), .A2(n6153), .ZN(n6356) );
  NAND2_X2 U3895 ( .A1(n6355), .A2(n6356), .ZN(n2478) );
  INV_X2 U3896 ( .A(n5062), .ZN(n6354) );
  NAND2_X2 U3902 ( .A1(n2478), .A2(n5066), .ZN(n827) );
  NAND2_X2 U3903 ( .A1(n3920), .A2(n1059), .ZN(n1286) );
  NOR2_X1 U3906 ( .A1(n3680), .A2(n4909), .ZN(n1467) );
  NOR2_X1 U3920 ( .A1(n1253), .A2(n2316), .ZN(n1249) );
  INV_X1 U3928 ( .A(n2316), .ZN(n1523) );
  BUF_X4 U3930 ( .A(n584), .Z(n6357) );
  NAND2_X2 U3932 ( .A1(n4913), .A2(n4914), .ZN(n1380) );
  INV_X2 U3933 ( .A(n4509), .ZN(n942) );
  INV_X2 U3934 ( .A(n4910), .ZN(n789) );
  NAND2_X2 U3935 ( .A1(n2120), .A2(n2119), .ZN(n2130) );
  NOR2_X2 U3938 ( .A1(n3653), .A2(n3652), .ZN(n3651) );
  NAND2_X4 U3939 ( .A1(n3179), .A2(n3182), .ZN(n3901) );
  OAI22_X1 U3940 ( .A1(n2622), .A2(n2623), .B1(n2621), .B2(n451), .ZN(n6358)
         );
  NAND2_X2 U3946 ( .A1(n3844), .A2(n3845), .ZN(n4278) );
  INV_X2 U3949 ( .A(n4298), .ZN(n4296) );
  INV_X2 U3960 ( .A(n5689), .ZN(n1008) );
  NAND2_X2 U3973 ( .A1(n4230), .A2(n4229), .ZN(n2971) );
  BUF_X2 U3992 ( .A(n5672), .Z(n6360) );
  NAND2_X2 U3995 ( .A1(n6361), .A2(n6362), .ZN(n6364) );
  NAND2_X2 U3998 ( .A1(n6363), .A2(n6364), .ZN(n4205) );
  INV_X1 U4015 ( .A(n1116), .ZN(n6362) );
  NAND2_X2 U4018 ( .A1(n4027), .A2(n2909), .ZN(n6365) );
  NOR2_X1 U4021 ( .A1(n3445), .A2(n566), .ZN(n3440) );
  INV_X1 U4039 ( .A(n3938), .ZN(n140) );
  INV_X2 U4042 ( .A(n5571), .ZN(n5862) );
  NAND2_X4 U4046 ( .A1(n122), .A2(n842), .ZN(n1548) );
  OR2_X2 U4048 ( .A1(n4473), .A2(n1754), .ZN(n989) );
  NAND2_X1 U4060 ( .A1(n2404), .A2(n5225), .ZN(n6369) );
  NAND2_X2 U4065 ( .A1(n6367), .A2(n6368), .ZN(n6370) );
  NAND2_X2 U4069 ( .A1(n6369), .A2(n6370), .ZN(n971) );
  INV_X2 U4080 ( .A(n2404), .ZN(n6367) );
  INV_X2 U4084 ( .A(n5332), .ZN(n2891) );
  INV_X1 U4096 ( .A(n2814), .ZN(n5370) );
  INV_X1 U4098 ( .A(n6609), .ZN(n2085) );
  NAND2_X1 U4102 ( .A1(n4339), .A2(n6609), .ZN(n2084) );
  OR2_X2 U4103 ( .A1(n4339), .A2(n3731), .ZN(n990) );
  NAND2_X1 U4135 ( .A1(n1771), .A2(n4117), .ZN(n6373) );
  INV_X1 U4154 ( .A(n4117), .ZN(n6372) );
  BUF_X4 U4158 ( .A(n5809), .Z(n6375) );
  NAND2_X2 U4162 ( .A1(n2941), .A2(n2940), .ZN(n6376) );
  NAND3_X1 U4164 ( .A1(n4099), .A2(b[0]), .A3(n397), .ZN(n1537) );
  NAND2_X2 U4168 ( .A1(n225), .A2(n226), .ZN(n6377) );
  NOR2_X2 U4175 ( .A1(n6093), .A2(n6092), .ZN(n5918) );
  NAND2_X1 U4191 ( .A1(n4735), .A2(n4736), .ZN(n561) );
  INV_X2 U4203 ( .A(n4735), .ZN(n559) );
  INV_X1 U4206 ( .A(n6332), .ZN(n6378) );
  NAND2_X2 U4207 ( .A1(n2298), .A2(n3983), .ZN(n6379) );
  NAND2_X2 U4209 ( .A1(n6432), .A2(n2470), .ZN(n6380) );
  BUF_X4 U4210 ( .A(n1915), .Z(n6381) );
  NAND2_X2 U4212 ( .A1(n4094), .A2(n6382), .ZN(n4101) );
  NOR2_X2 U4249 ( .A1(n6384), .A2(n6383), .ZN(n6382) );
  NOR2_X2 U4265 ( .A1(n4405), .A2(n3538), .ZN(n6384) );
  NAND2_X2 U4270 ( .A1(n2652), .A2(n4451), .ZN(n6385) );
  NAND2_X2 U4272 ( .A1(n6386), .A2(n1584), .ZN(n1087) );
  NAND2_X2 U4289 ( .A1(n2852), .A2(n1485), .ZN(n2422) );
  NAND2_X2 U4291 ( .A1(n5037), .A2(n5038), .ZN(n2852) );
  NAND2_X2 U4301 ( .A1(n6388), .A2(n6387), .ZN(n4173) );
  NAND2_X2 U4319 ( .A1(n4506), .A2(b[3]), .ZN(n6388) );
  NAND2_X2 U4331 ( .A1(n6390), .A2(n2027), .ZN(n4730) );
  NAND3_X2 U4339 ( .A1(n1705), .A2(n1703), .A3(n1704), .ZN(n2026) );
  BUF_X4 U4340 ( .A(n3608), .Z(n6391) );
  NAND2_X1 U4341 ( .A1(n4633), .A2(n4632), .ZN(n1990) );
  NAND2_X2 U4343 ( .A1(n3339), .A2(n3336), .ZN(n4633) );
  NOR3_X4 U4353 ( .A1(n3298), .A2(a[16]), .A3(a[15]), .ZN(n4768) );
  NAND2_X2 U4354 ( .A1(n6392), .A2(n443), .ZN(n1199) );
  NAND2_X2 U4367 ( .A1(n2792), .A2(n4564), .ZN(n6392) );
  NOR2_X2 U4369 ( .A1(n4947), .A2(n6393), .ZN(n3088) );
  NOR2_X2 U4382 ( .A1(n5190), .A2(n4945), .ZN(n6393) );
  NAND2_X2 U4400 ( .A1(n1466), .A2(n4686), .ZN(n3550) );
  NOR3_X2 U4419 ( .A1(n5089), .A2(n5088), .A3(n258), .ZN(n2797) );
  NAND2_X4 U4430 ( .A1(n2179), .A2(n2178), .ZN(n1278) );
  NAND2_X4 U4432 ( .A1(n1563), .A2(n6394), .ZN(n1870) );
  INV_X4 U4435 ( .A(n1817), .ZN(n6394) );
  NOR2_X2 U4443 ( .A1(n1789), .A2(n1131), .ZN(n1817) );
  INV_X4 U4445 ( .A(n6395), .ZN(n2683) );
  NOR2_X2 U4454 ( .A1(n3222), .A2(n4711), .ZN(n6395) );
  NAND2_X2 U4463 ( .A1(n1472), .A2(n1471), .ZN(n3222) );
  NAND2_X2 U4475 ( .A1(n6397), .A2(n6163), .ZN(n1826) );
  NAND2_X2 U4480 ( .A1(n1207), .A2(n4705), .ZN(n6397) );
  AOI21_X2 U4496 ( .B1(n4275), .B2(n4276), .A(n4274), .ZN(n4282) );
  NOR2_X2 U4508 ( .A1(n1507), .A2(n1627), .ZN(n6398) );
  NAND2_X2 U4516 ( .A1(n2046), .A2(n2047), .ZN(n6399) );
  NAND3_X2 U4535 ( .A1(n2136), .A2(n2134), .A3(n2137), .ZN(n2429) );
  NAND2_X4 U4540 ( .A1(n6401), .A2(n6400), .ZN(n4368) );
  INV_X2 U4553 ( .A(n4360), .ZN(n6400) );
  NAND2_X2 U4561 ( .A1(n4361), .A2(a[0]), .ZN(n6401) );
  INV_X2 U4569 ( .A(n1658), .ZN(n567) );
  NOR2_X2 U4575 ( .A1(n4804), .A2(n3103), .ZN(n1757) );
  OAI21_X2 U4589 ( .B1(n2924), .B2(n4490), .A(n2923), .ZN(n4453) );
  AOI22_X2 U4594 ( .A1(n1386), .A2(n4663), .B1(n1438), .B2(n1387), .ZN(n2773)
         );
  NAND2_X2 U4602 ( .A1(n856), .A2(n855), .ZN(n4298) );
  NOR2_X2 U4604 ( .A1(n2114), .A2(n4280), .ZN(n4299) );
  NAND2_X2 U4607 ( .A1(n2177), .A2(n1278), .ZN(n2174) );
  AOI21_X2 U4628 ( .B1(n1976), .B2(n4627), .A(n97), .ZN(n2535) );
  NAND2_X2 U4675 ( .A1(n6607), .A2(n2150), .ZN(n1334) );
  NOR2_X2 U4690 ( .A1(n1078), .A2(n1077), .ZN(n6405) );
  NAND2_X2 U4693 ( .A1(n1926), .A2(n2470), .ZN(n142) );
  NAND2_X2 U4697 ( .A1(n3254), .A2(n148), .ZN(n1926) );
  NAND2_X2 U4698 ( .A1(n1061), .A2(n3513), .ZN(n2336) );
  NOR2_X4 U4736 ( .A1(n2337), .A2(n4812), .ZN(n3513) );
  NAND2_X2 U4749 ( .A1(n4244), .A2(n4308), .ZN(n3034) );
  BUF_X4 U4759 ( .A(n4724), .Z(n6406) );
  NAND2_X2 U4760 ( .A1(n3127), .A2(n4761), .ZN(n6407) );
  OAI21_X2 U4789 ( .B1(n3386), .B2(n4741), .A(n3469), .ZN(n1987) );
  NAND2_X1 U4803 ( .A1(n5260), .A2(n5259), .ZN(n456) );
  NAND2_X2 U4807 ( .A1(n6408), .A2(n2385), .ZN(n2575) );
  NAND2_X2 U4808 ( .A1(n4078), .A2(n1115), .ZN(n6408) );
  NAND3_X2 U4901 ( .A1(n6410), .A2(n2690), .A3(n2691), .ZN(n1601) );
  INV_X4 U4903 ( .A(n4528), .ZN(n6410) );
  NAND2_X4 U4910 ( .A1(n2040), .A2(n2039), .ZN(n4528) );
  NOR3_X4 U4923 ( .A1(n6411), .A2(n187), .A3(a[13]), .ZN(n3022) );
  INV_X4 U4931 ( .A(a[11]), .ZN(n6411) );
  NAND2_X2 U4932 ( .A1(n4939), .A2(n4938), .ZN(n1758) );
  OAI22_X2 U4941 ( .A1(n4809), .A2(n341), .B1(n4807), .B2(n139), .ZN(n4938) );
  INV_X2 U4948 ( .A(n6412), .ZN(n439) );
  NAND2_X2 U4958 ( .A1(n3831), .A2(n3833), .ZN(n6412) );
  NOR2_X2 U4963 ( .A1(n2132), .A2(n2139), .ZN(n2428) );
  AOI21_X2 U4966 ( .B1(n2140), .B2(n3462), .A(n4273), .ZN(n2139) );
  NOR2_X2 U4969 ( .A1(n4445), .A2(n3604), .ZN(n3349) );
  BUF_X4 U4978 ( .A(n5374), .Z(n6413) );
  NOR2_X2 U4985 ( .A1(n5360), .A2(n4794), .ZN(n6415) );
  NAND3_X2 U4998 ( .A1(n3976), .A2(n793), .A3(n792), .ZN(n615) );
  AOI21_X2 U4999 ( .B1(n3838), .B2(n3764), .A(n4271), .ZN(n3463) );
  NOR2_X2 U5003 ( .A1(n3836), .A2(n3837), .ZN(n3838) );
  NAND2_X2 U5004 ( .A1(n6530), .A2(n534), .ZN(n537) );
  INV_X2 U5028 ( .A(n6417), .ZN(n3138) );
  NAND2_X2 U5043 ( .A1(n1145), .A2(n4970), .ZN(n6417) );
  NAND2_X2 U5051 ( .A1(n2731), .A2(n1059), .ZN(n6418) );
  NAND2_X2 U5054 ( .A1(n6419), .A2(n889), .ZN(n5251) );
  NAND2_X2 U5068 ( .A1(n887), .A2(n888), .ZN(n6419) );
  NAND2_X2 U5071 ( .A1(n6420), .A2(n5185), .ZN(n5246) );
  NOR2_X2 U5073 ( .A1(n2204), .A2(n2203), .ZN(n6420) );
  NOR2_X2 U5074 ( .A1(n6421), .A2(n2346), .ZN(n3509) );
  NOR2_X2 U5075 ( .A1(n239), .A2(n4377), .ZN(n6421) );
  INV_X4 U5076 ( .A(n6422), .ZN(n1948) );
  NOR2_X2 U5077 ( .A1(n3319), .A2(n2852), .ZN(n6422) );
  NAND2_X2 U5079 ( .A1(n3550), .A2(n707), .ZN(n4903) );
  NAND2_X2 U5095 ( .A1(n1952), .A2(n1951), .ZN(n2613) );
  BUF_X4 U5100 ( .A(n6325), .Z(n6423) );
  OR2_X2 U5111 ( .A1(n5219), .A2(b[18]), .ZN(n1392) );
  BUF_X4 U5119 ( .A(n5255), .Z(n6424) );
  NOR2_X2 U5121 ( .A1(n1395), .A2(n6425), .ZN(n5187) );
  NAND2_X2 U5122 ( .A1(n6427), .A2(n6426), .ZN(n6425) );
  NAND2_X2 U5130 ( .A1(n2537), .A2(b[15]), .ZN(n6426) );
  OAI21_X2 U5135 ( .B1(n4589), .B2(n1529), .A(n3711), .ZN(n6432) );
  NOR2_X4 U5140 ( .A1(n1527), .A2(n1528), .ZN(n4589) );
  NAND2_X2 U5148 ( .A1(n6465), .A2(n6428), .ZN(n232) );
  INV_X2 U5165 ( .A(n4670), .ZN(n6428) );
  NOR2_X2 U5168 ( .A1(n2441), .A2(n1428), .ZN(n1889) );
  NAND2_X2 U5172 ( .A1(n5139), .A2(n5138), .ZN(n2441) );
  NAND2_X2 U5185 ( .A1(n1510), .A2(n1509), .ZN(n3640) );
  NAND2_X2 U5195 ( .A1(n2232), .A2(n2886), .ZN(n1510) );
  INV_X2 U5202 ( .A(n1935), .ZN(n943) );
  OAI21_X2 U5205 ( .B1(n4396), .B2(n4395), .A(n3327), .ZN(n1935) );
  INV_X2 U5207 ( .A(n5259), .ZN(n6431) );
  OAI21_X2 U5211 ( .B1(n3181), .B2(n2980), .A(n2979), .ZN(n4686) );
  NAND2_X2 U5213 ( .A1(n6433), .A2(n316), .ZN(n318) );
  INV_X2 U5225 ( .A(n1565), .ZN(n6433) );
  INV_X2 U5255 ( .A(n6434), .ZN(n1683) );
  NAND2_X2 U5261 ( .A1(n4905), .A2(n4906), .ZN(n6434) );
  NAND2_X2 U5272 ( .A1(n6435), .A2(n3561), .ZN(n1156) );
  NAND2_X2 U5275 ( .A1(n88), .A2(n2090), .ZN(n6435) );
  OAI21_X2 U5279 ( .B1(n2091), .B2(n3015), .A(n2131), .ZN(n2090) );
  NAND2_X2 U5283 ( .A1(n711), .A2(n4475), .ZN(n6437) );
  NAND2_X2 U5294 ( .A1(n2591), .A2(n2592), .ZN(n6438) );
  BUF_X4 U5295 ( .A(n4887), .Z(n6439) );
  NAND2_X2 U5335 ( .A1(n1709), .A2(n2901), .ZN(n6442) );
  INV_X2 U5376 ( .A(n2074), .ZN(n6443) );
  NOR3_X2 U5377 ( .A1(n3667), .A2(n3668), .A3(n3435), .ZN(n3666) );
  INV_X4 U5378 ( .A(b[20]), .ZN(n5471) );
  MUX2_X2 U5396 ( .A(n512), .B(n606), .S(b[20]), .Z(n4771) );
  OAI22_X2 U5405 ( .A1(n6444), .A2(n4490), .B1(n471), .B2(b[20]), .ZN(n4329)
         );
  XNOR2_X2 U5406 ( .A(a[1]), .B(b[21]), .ZN(n6444) );
  NOR2_X2 U5407 ( .A1(a[1]), .A2(a[2]), .ZN(n1358) );
  INV_X2 U5408 ( .A(n1689), .ZN(n154) );
  XOR2_X2 U5435 ( .A(a[11]), .B(b[4]), .Z(n6445) );
  INV_X4 U5453 ( .A(n4073), .ZN(n818) );
  NOR2_X4 U5462 ( .A1(n5101), .A2(a[11]), .ZN(n440) );
  INV_X2 U5472 ( .A(n5246), .ZN(n888) );
  INV_X1 U5481 ( .A(n5265), .ZN(n2499) );
  AND2_X4 U5483 ( .A1(n2938), .A2(n2937), .ZN(n6447) );
  INV_X4 U5509 ( .A(n3260), .ZN(n3013) );
  INV_X2 U5544 ( .A(n4871), .ZN(n689) );
  INV_X4 U5545 ( .A(n5561), .ZN(n5558) );
  INV_X4 U5547 ( .A(n5330), .ZN(n660) );
  OR2_X2 U5587 ( .A1(n5090), .A2(n5089), .ZN(n6451) );
  AND2_X2 U5591 ( .A1(n5029), .A2(n2751), .ZN(n6452) );
  INV_X2 U5597 ( .A(n1954), .ZN(n3075) );
  INV_X4 U5619 ( .A(n3930), .ZN(n762) );
  INV_X4 U5621 ( .A(n5130), .ZN(n280) );
  AOI21_X2 U5622 ( .B1(n5176), .B2(n5177), .A(n3384), .ZN(n639) );
  INV_X4 U5625 ( .A(n4968), .ZN(n690) );
  NAND2_X4 U5628 ( .A1(n3467), .A2(n1470), .ZN(n2003) );
  INV_X2 U5633 ( .A(n5839), .ZN(n1015) );
  NAND2_X2 U5634 ( .A1(n3269), .A2(n5030), .ZN(n3748) );
  NOR2_X4 U5636 ( .A1(n1262), .A2(n1263), .ZN(n3200) );
  INV_X1 U5638 ( .A(n2154), .ZN(n2155) );
  NOR2_X4 U5655 ( .A1(n1548), .A2(n4313), .ZN(n5707) );
  NAND2_X2 U3490 ( .A1(n984), .A2(n4940), .ZN(n4849) );
  NOR2_X4 U3272 ( .A1(n1275), .A2(n2223), .ZN(n4377) );
  OAI21_X2 U1076 ( .B1(n4377), .B2(n4376), .A(n4375), .ZN(n4474) );
  NAND2_X4 U4877 ( .A1(n564), .A2(n4431), .ZN(n4432) );
  INV_X4 U2235 ( .A(n4388), .ZN(n1833) );
  NOR2_X2 U4929 ( .A1(n4434), .A2(n3598), .ZN(n2776) );
  NAND2_X2 U1450 ( .A1(n2697), .A2(n6621), .ZN(n6215) );
  INV_X8 U677 ( .A(n817), .ZN(n564) );
  NOR2_X4 U1019 ( .A1(n4521), .A2(n458), .ZN(n1184) );
  INV_X4 U2942 ( .A(n5085), .ZN(n6303) );
  NAND2_X4 U2164 ( .A1(n207), .A2(n833), .ZN(n835) );
  NAND2_X4 U1130 ( .A1(n5599), .A2(n5597), .ZN(n5927) );
  OAI22_X2 U5575 ( .A1(n5205), .A2(n5204), .B1(n5203), .B2(n1103), .ZN(n5207)
         );
  NAND2_X2 U1991 ( .A1(n5042), .A2(n3632), .ZN(n686) );
  INV_X4 U3574 ( .A(n2244), .ZN(n47) );
  NAND2_X2 U1987 ( .A1(n5077), .A2(b[16]), .ZN(n3401) );
  NAND2_X2 U1593 ( .A1(n2318), .A2(n4523), .ZN(n2107) );
  AOI22_X2 U3641 ( .A1(n3835), .A2(n3230), .B1(b[5]), .B2(n5136), .ZN(n2801)
         );
  INV_X4 U708 ( .A(n4912), .ZN(n138) );
  INV_X4 U1051 ( .A(n1894), .ZN(n1953) );
  INV_X2 U2112 ( .A(n4579), .ZN(n2610) );
  INV_X2 U1841 ( .A(n2323), .ZN(n939) );
  NAND2_X2 U1510 ( .A1(n1688), .A2(n4269), .ZN(n3033) );
  NOR2_X4 U1895 ( .A1(n3923), .A2(n3922), .ZN(n6251) );
  NOR2_X4 U4565 ( .A1(n4668), .A2(n1696), .ZN(n2536) );
  NAND2_X2 U2477 ( .A1(n1666), .A2(n1665), .ZN(n6288) );
  NAND2_X4 U1115 ( .A1(n2457), .A2(n2456), .ZN(n3152) );
  NAND2_X4 U3112 ( .A1(n4688), .A2(n3562), .ZN(n1163) );
  NAND2_X2 U1779 ( .A1(n1070), .A2(n1069), .ZN(n590) );
  NOR2_X4 U2376 ( .A1(n3598), .A2(n4548), .ZN(n2467) );
  NOR3_X4 U1414 ( .A1(n1248), .A2(a[1]), .A3(a[2]), .ZN(n568) );
  NOR2_X4 U24 ( .A1(n365), .A2(a[3]), .ZN(n6211) );
  NAND2_X4 U4093 ( .A1(n1449), .A2(n30), .ZN(n2001) );
  NOR2_X2 U2739 ( .A1(n4969), .A2(n1089), .ZN(n5805) );
  NOR2_X4 U4568 ( .A1(n5266), .A2(b[6]), .ZN(n2622) );
  NAND2_X4 U2506 ( .A1(n3094), .A2(n4024), .ZN(n4451) );
  NOR2_X4 U1253 ( .A1(n3808), .A2(n3807), .ZN(n1865) );
  INV_X4 U3253 ( .A(n1651), .ZN(n1261) );
  INV_X4 U2968 ( .A(n4328), .ZN(n6304) );
  INV_X4 U2328 ( .A(n1125), .ZN(n904) );
  XOR2_X2 U1348 ( .A(n4883), .B(n1440), .Z(n6204) );
  NOR2_X4 U4094 ( .A1(n5859), .A2(n5860), .ZN(n5854) );
  NAND2_X2 U1873 ( .A1(n3483), .A2(n5548), .ZN(n623) );
  OAI21_X2 U4726 ( .B1(n4117), .B2(n4116), .A(n4114), .ZN(n4113) );
  NAND2_X4 U764 ( .A1(n399), .A2(n1766), .ZN(n4191) );
  NOR2_X4 U4613 ( .A1(n5366), .A2(n5365), .ZN(n5458) );
  OAI21_X2 U1881 ( .B1(n5550), .B2(n5549), .A(n966), .ZN(n5548) );
  NAND2_X2 U5044 ( .A1(n5385), .A2(n680), .ZN(n5393) );
  NAND2_X2 U1985 ( .A1(n6492), .A2(n5808), .ZN(n680) );
  NAND2_X2 U4662 ( .A1(n4507), .A2(n6528), .ZN(n4511) );
  NOR2_X2 U1868 ( .A1(n5493), .A2(n5492), .ZN(n5550) );
  NOR2_X2 U1838 ( .A1(n3699), .A2(n5267), .ZN(n5268) );
  INV_X4 U4214 ( .A(n6092), .ZN(n2156) );
  NAND2_X2 U1525 ( .A1(n4238), .A2(b[13]), .ZN(n1737) );
  INV_X4 U3884 ( .A(n3912), .ZN(n1056) );
  OAI21_X2 U4775 ( .B1(n4658), .B2(n5105), .A(n4661), .ZN(n4660) );
  NOR2_X2 U5269 ( .A1(n3431), .A2(b[19]), .ZN(n3436) );
  NAND3_X2 U1030 ( .A1(n4167), .A2(n4165), .A3(n4166), .ZN(n4171) );
  NAND2_X2 U4131 ( .A1(n4163), .A2(n4164), .ZN(n4167) );
  INV_X4 U4467 ( .A(n2855), .ZN(n2485) );
  NAND3_X2 U1520 ( .A1(n818), .A2(n1294), .A3(n1295), .ZN(n6227) );
  INV_X4 U1210 ( .A(n4322), .ZN(n291) );
  INV_X4 U1049 ( .A(n3083), .ZN(n2901) );
  NAND2_X4 U1129 ( .A1(n5599), .A2(n5597), .ZN(n259) );
  NOR2_X2 U4481 ( .A1(n1058), .A2(n2602), .ZN(n2509) );
  INV_X4 U136 ( .A(n4872), .ZN(n913) );
  INV_X4 U1474 ( .A(n4108), .ZN(n426) );
  NOR2_X2 U1572 ( .A1(n513), .A2(n4794), .ZN(n4931) );
  NAND2_X2 U2356 ( .A1(n1230), .A2(n461), .ZN(n933) );
  INV_X2 U1753 ( .A(n1628), .ZN(n570) );
  INV_X4 U1309 ( .A(n4038), .ZN(n334) );
  NAND2_X2 U3046 ( .A1(n1194), .A2(b[12]), .ZN(n1111) );
  NAND2_X2 U2444 ( .A1(n4840), .A2(n973), .ZN(n4792) );
  NAND2_X2 U1221 ( .A1(n1662), .A2(n4926), .ZN(n302) );
  NOR2_X4 U4012 ( .A1(n2056), .A2(n2256), .ZN(n2549) );
  INV_X4 U113 ( .A(n5507), .ZN(n5505) );
  INV_X4 U1874 ( .A(n3483), .ZN(n621) );
  NAND2_X4 U5399 ( .A1(n5546), .A2(n5547), .ZN(n3483) );
  NAND2_X4 U1502 ( .A1(n1915), .A2(n5662), .ZN(n5667) );
  INV_X4 U2358 ( .A(n1230), .ZN(n932) );
  INV_X4 U4148 ( .A(n2059), .ZN(n2338) );
  INV_X4 U1428 ( .A(n2826), .ZN(n6214) );
  NAND2_X4 U1260 ( .A1(n4689), .A2(n4389), .ZN(n4045) );
  INV_X8 U1085 ( .A(n2854), .ZN(n2829) );
  NAND2_X2 U5035 ( .A1(n639), .A2(n6192), .ZN(n5261) );
  NOR2_X4 U2753 ( .A1(n1005), .A2(n1009), .ZN(n4670) );
  OAI21_X2 U369 ( .B1(n2481), .B2(n3546), .A(n1005), .ZN(n6287) );
  INV_X8 U2201 ( .A(n3152), .ZN(n1009) );
  NOR2_X4 U557 ( .A1(n2950), .A2(n1324), .ZN(n2623) );
  OAI22_X2 U4755 ( .A1(n4676), .A2(n4675), .B1(n4835), .B2(n6406), .ZN(n4683)
         );
  NOR2_X4 U1511 ( .A1(a[11]), .A2(n360), .ZN(n2675) );
  NAND2_X2 U2012 ( .A1(n4303), .A2(n1026), .ZN(n901) );
  NAND2_X4 U2387 ( .A1(n3470), .A2(n4728), .ZN(n3250) );
  NAND2_X2 U4398 ( .A1(n880), .A2(n879), .ZN(n1465) );
  NAND2_X4 U1052 ( .A1(n665), .A2(n664), .ZN(n1894) );
  NOR2_X4 U5438 ( .A1(n2656), .A2(b[1]), .ZN(n3544) );
  INV_X4 U354 ( .A(n3229), .ZN(n2896) );
  INV_X4 U582 ( .A(n2803), .ZN(n3171) );
  NAND2_X4 U1107 ( .A1(n250), .A2(n364), .ZN(n3229) );
  INV_X4 U3211 ( .A(n2350), .ZN(n4839) );
  NAND2_X4 U652 ( .A1(n1898), .A2(n1897), .ZN(n1628) );
  NAND2_X2 U1178 ( .A1(n4908), .A2(n4907), .ZN(n1897) );
  INV_X4 U140 ( .A(n1222), .ZN(n518) );
  XNOR2_X2 U2823 ( .A(n1628), .B(n4916), .ZN(n2447) );
  NAND2_X2 U1672 ( .A1(n1222), .A2(n4867), .ZN(n520) );
  NOR2_X2 U391 ( .A1(b[3]), .A2(n6326), .ZN(n4421) );
  NOR2_X2 U190 ( .A1(n4635), .A2(n4637), .ZN(n4480) );
  NAND2_X4 U3387 ( .A1(n5735), .A2(n5733), .ZN(n6325) );
  NAND2_X2 U1231 ( .A1(n792), .A2(n793), .ZN(n304) );
  OAI21_X2 U4741 ( .B1(n5845), .B2(n1099), .A(n5844), .ZN(n5846) );
  NOR3_X2 U1685 ( .A1(n2772), .A2(n4665), .A3(n3152), .ZN(n2771) );
  INV_X8 U97 ( .A(b[12]), .ZN(n5277) );
  INV_X4 U2827 ( .A(n4516), .ZN(n4518) );
  INV_X2 U1323 ( .A(n3655), .ZN(n1913) );
  INV_X2 U5201 ( .A(n3322), .ZN(n3123) );
  NAND2_X2 U2167 ( .A1(n1566), .A2(n4466), .ZN(n797) );
  NAND2_X4 U4174 ( .A1(n151), .A2(n848), .ZN(n226) );
  OAI21_X2 U2403 ( .B1(n3579), .B2(n891), .A(n3578), .ZN(n5093) );
  INV_X4 U1763 ( .A(n3604), .ZN(n577) );
  INV_X4 U4267 ( .A(n4444), .ZN(n2220) );
  NOR2_X4 U2752 ( .A1(n3331), .A2(n3256), .ZN(n3332) );
  NOR2_X4 U2791 ( .A1(n2987), .A2(n2373), .ZN(n3322) );
  NAND2_X2 U2368 ( .A1(n4687), .A2(a[13]), .ZN(n4364) );
  NOR2_X2 U4750 ( .A1(n760), .A2(n3538), .ZN(n4420) );
  NOR2_X2 U1930 ( .A1(n4060), .A2(n4059), .ZN(n4058) );
  INV_X8 U4683 ( .A(n4795), .ZN(n4746) );
  NOR3_X2 U4661 ( .A1(a[0]), .A2(b[19]), .A3(n2695), .ZN(n4360) );
  NAND2_X4 U1694 ( .A1(n798), .A2(n797), .ZN(n1843) );
  NAND2_X4 U2171 ( .A1(n4810), .A2(b[12]), .ZN(n4347) );
  INV_X4 U226 ( .A(n4371), .ZN(n4370) );
  NOR2_X4 U922 ( .A1(n1843), .A2(n1842), .ZN(n1841) );
  NAND2_X2 U5288 ( .A1(n2715), .A2(n1059), .ZN(n3225) );
  NAND2_X4 U49 ( .A1(n397), .A2(n6162), .ZN(n399) );
  NAND2_X2 U1660 ( .A1(n5295), .A2(n5294), .ZN(n1732) );
  INV_X4 U2000 ( .A(n1945), .ZN(n3726) );
  NAND2_X2 U17 ( .A1(a[23]), .A2(b[20]), .ZN(n5957) );
  INV_X4 U1244 ( .A(a[15]), .ZN(n310) );
  NAND2_X1 U2917 ( .A1(b[19]), .A2(b[18]), .ZN(n5905) );
  INV_X1 U334 ( .A(b[15]), .ZN(n35) );
  NAND2_X1 U2524 ( .A1(b[13]), .A2(b[12]), .ZN(n5344) );
  OAI21_X1 U2904 ( .B1(b[12]), .B2(b[13]), .A(a[23]), .ZN(n5343) );
  NAND2_X1 U2396 ( .A1(b[15]), .A2(b[14]), .ZN(n5470) );
  NAND2_X2 U3652 ( .A1(n6340), .A2(n6341), .ZN(n6343) );
  INV_X2 U2017 ( .A(n3258), .ZN(n704) );
  NAND2_X2 U1645 ( .A1(a[14]), .A2(n502), .ZN(n503) );
  AND2_X2 U1147 ( .A1(n6182), .A2(a[7]), .ZN(n267) );
  AND2_X2 U2458 ( .A1(n267), .A2(n4942), .ZN(n988) );
  OR2_X2 U2414 ( .A1(n465), .A2(n3572), .ZN(n946) );
  INV_X4 U3100 ( .A(n3022), .ZN(n1147) );
  NAND2_X2 U1243 ( .A1(n312), .A2(n313), .ZN(n3507) );
  INV_X2 U3316 ( .A(n2675), .ZN(n6322) );
  INV_X2 U1575 ( .A(n6415), .ZN(n6231) );
  NOR2_X2 U2025 ( .A1(n4502), .A2(n4501), .ZN(n2486) );
  INV_X2 U3200 ( .A(n4854), .ZN(n1220) );
  AND2_X2 U715 ( .A1(n6242), .A2(n6528), .ZN(n6157) );
  OR2_X2 U4884 ( .A1(n3631), .A2(n3630), .ZN(n2703) );
  INV_X2 U2842 ( .A(n4214), .ZN(n4215) );
  NAND3_X2 U3678 ( .A1(n3841), .A2(n2746), .A3(n2142), .ZN(n4273) );
  INV_X2 U559 ( .A(n2792), .ZN(n1280) );
  INV_X2 U1171 ( .A(n1045), .ZN(n282) );
  INV_X4 U1099 ( .A(n4760), .ZN(n245) );
  INV_X2 U3471 ( .A(n4273), .ZN(n3464) );
  NAND2_X2 U958 ( .A1(n1192), .A2(n1191), .ZN(n2503) );
  NAND2_X1 U6164 ( .A1(n195), .A2(n6034), .ZN(n6047) );
  NOR2_X2 U2927 ( .A1(n6414), .A2(n4827), .ZN(n4874) );
  INV_X2 U2820 ( .A(n4404), .ZN(n3693) );
  INV_X2 U4913 ( .A(n5025), .ZN(n2753) );
  INV_X2 U3357 ( .A(n2432), .ZN(n1549) );
  NOR2_X2 U2298 ( .A1(n2464), .A2(n2463), .ZN(n4652) );
  NAND2_X2 U1628 ( .A1(n5271), .A2(n5270), .ZN(n5351) );
  INV_X2 U753 ( .A(n2634), .ZN(n6167) );
  NAND2_X2 U762 ( .A1(n6167), .A2(n4864), .ZN(n1558) );
  INV_X2 U2216 ( .A(n5066), .ZN(n826) );
  XNOR2_X1 U2772 ( .A(n6106), .B(n6105), .ZN(n6124) );
  NAND2_X2 U4945 ( .A1(n4804), .A2(n3103), .ZN(n4939) );
  NAND2_X2 U3415 ( .A1(n429), .A2(n428), .ZN(n1540) );
  INV_X2 U401 ( .A(n4374), .ZN(n2907) );
  NAND2_X2 U1506 ( .A1(n819), .A2(n6227), .ZN(n1367) );
  NAND2_X2 U3942 ( .A1(n3844), .A2(n3845), .ZN(n6359) );
  NOR2_X1 U2734 ( .A1(n5940), .A2(n5943), .ZN(n5946) );
  NOR2_X2 U236 ( .A1(n1583), .A2(n3064), .ZN(n1484) );
  NOR2_X2 U853 ( .A1(n1367), .A2(n2636), .ZN(n177) );
  BUF_X2 U201 ( .A(n5202), .Z(n1103) );
  AOI21_X1 U698 ( .B1(n6117), .B2(n6052), .A(n6116), .ZN(n6053) );
  AND2_X2 U4860 ( .A1(n6108), .A2(n6051), .ZN(n6049) );
  OR2_X2 U154 ( .A1(n3948), .A2(n3746), .ZN(n991) );
  INV_X2 U1875 ( .A(n5548), .ZN(n622) );
  NAND2_X2 U156 ( .A1(n2969), .A2(n2968), .ZN(n1845) );
  INV_X2 U3052 ( .A(n2387), .ZN(n1115) );
  INV_X2 U3980 ( .A(n4643), .ZN(n2164) );
  NAND2_X2 U3175 ( .A1(n1654), .A2(n2765), .ZN(n1202) );
  INV_X2 U5505 ( .A(n5563), .ZN(n3191) );
  INV_X2 U1212 ( .A(n5547), .ZN(n5515) );
  INV_X2 U1587 ( .A(n6257), .ZN(n969) );
  AOI21_X1 U5827 ( .B1(n4647), .B2(n6604), .A(n4645), .ZN(n4648) );
  INV_X2 U2005 ( .A(n1665), .ZN(n692) );
  XNOR2_X1 U2679 ( .A(n3590), .B(n64), .ZN(n5736) );
  INV_X1 U2686 ( .A(n3167), .ZN(n5712) );
  NAND2_X1 U4614 ( .A1(n5730), .A2(n6423), .ZN(n5731) );
  XNOR2_X2 U5432 ( .A(n6491), .B(n1085), .ZN(n5812) );
  INV_X2 U4739 ( .A(n5812), .ZN(n3140) );
  NAND2_X2 U5137 ( .A1(n6661), .A2(n736), .ZN(n5627) );
  INV_X1 U2353 ( .A(n5373), .ZN(n926) );
  INV_X2 U5897 ( .A(n6613), .ZN(n5853) );
  XNOR2_X1 U4851 ( .A(n5615), .B(n5616), .ZN(n5613) );
  INV_X2 U4742 ( .A(n5843), .ZN(n5844) );
  INV_X2 U4922 ( .A(n2864), .ZN(n5924) );
  AND2_X1 U383 ( .A1(n1013), .A2(n6661), .ZN(n2728) );
  NAND2_X2 U5528 ( .A1(n2745), .A2(n6459), .ZN(n3739) );
  NOR2_X4 U4292 ( .A1(n6436), .A2(n4476), .ZN(n1154) );
  XNOR2_X2 U3627 ( .A(n4616), .B(n4544), .ZN(n2147) );
  INV_X4 U953 ( .A(n1747), .ZN(n207) );
  INV_X4 U891 ( .A(n3619), .ZN(n2112) );
  NAND2_X4 U8 ( .A1(n1269), .A2(n6222), .ZN(n3382) );
  INV_X4 U1557 ( .A(a[11]), .ZN(n3826) );
  INV_X4 U5428 ( .A(b[18]), .ZN(n5529) );
  INV_X4 U3518 ( .A(n1405), .ZN(n4812) );
  NAND2_X2 U1242 ( .A1(n310), .A2(a[16]), .ZN(n313) );
  NAND2_X2 U5589 ( .A1(a[1]), .A2(a[2]), .ZN(n4021) );
  NAND2_X2 U5256 ( .A1(n4026), .A2(a[17]), .ZN(n4424) );
  NOR2_X2 U148 ( .A1(n4674), .A2(a[3]), .ZN(n4678) );
  NAND2_X2 U5590 ( .A1(n4021), .A2(n4492), .ZN(n3773) );
  NAND2_X2 U86 ( .A1(n3507), .A2(a[17]), .ZN(n314) );
  NAND2_X2 U5867 ( .A1(n5951), .A2(a[7]), .ZN(n4817) );
  INV_X4 U494 ( .A(n4600), .ZN(n6155) );
  NOR2_X2 U2969 ( .A1(n267), .A2(b[20]), .ZN(n4741) );
  NAND2_X2 U5959 ( .A1(n5232), .A2(n5231), .ZN(n5284) );
  NOR2_X2 U862 ( .A1(n2602), .A2(b[1]), .ZN(n2507) );
  NOR2_X2 U60 ( .A1(n2656), .A2(b[12]), .ZN(n2400) );
  NAND2_X2 U1872 ( .A1(n5900), .A2(b[1]), .ZN(n3086) );
  NOR2_X2 U3614 ( .A1(n2507), .A2(n4189), .ZN(n2506) );
  NOR2_X2 U43 ( .A1(n2995), .A2(n1717), .ZN(n3380) );
  NOR2_X2 U1862 ( .A1(n6251), .A2(n3965), .ZN(n1969) );
  NAND2_X2 U3297 ( .A1(n1292), .A2(n1290), .ZN(n4073) );
  NOR2_X2 U2147 ( .A1(n4103), .A2(n4104), .ZN(n4108) );
  NAND2_X2 U36 ( .A1(n1139), .A2(n2509), .ZN(n4231) );
  NAND2_X2 U170 ( .A1(n4433), .A2(n4432), .ZN(n4449) );
  NOR2_X2 U135 ( .A1(n5505), .A2(n5504), .ZN(n5552) );
  NOR2_X2 U5931 ( .A1(n1032), .A2(n5121), .ZN(n5125) );
  NAND2_X2 U682 ( .A1(n1025), .A2(n3410), .ZN(n1240) );
  NAND2_X2 U2159 ( .A1(n835), .A2(n834), .ZN(n1374) );
  NAND2_X2 U805 ( .A1(n5580), .A2(n5581), .ZN(n6000) );
  NOR2_X2 U3271 ( .A1(n1274), .A2(n3553), .ZN(n5375) );
  NOR2_X2 U1411 ( .A1(n5808), .A2(n3391), .ZN(n2783) );
  NAND2_X2 U9 ( .A1(n3690), .A2(n5083), .ZN(n5084) );
  NAND2_X2 U14 ( .A1(n3052), .A2(n3058), .ZN(n2606) );
  NAND3_X2 U16 ( .A1(n1916), .A2(a[12]), .A3(a[11]), .ZN(n4774) );
  NAND2_X2 U20 ( .A1(a[7]), .A2(n6606), .ZN(n6605) );
  INV_X4 U31 ( .A(b[17]), .ZN(n6515) );
  INV_X4 U32 ( .A(a[10]), .ZN(n466) );
  INV_X4 U42 ( .A(a[12]), .ZN(n2684) );
  NAND3_X2 U47 ( .A1(n256), .A2(n6525), .A3(n3759), .ZN(n152) );
  NAND2_X4 U56 ( .A1(n3926), .A2(n6593), .ZN(n3940) );
  XNOR2_X2 U62 ( .A(n5687), .B(n5686), .ZN(\d[10]_BAR ) );
  NOR2_X2 U66 ( .A1(n365), .A2(a[3]), .ZN(n648) );
  AND2_X4 U67 ( .A1(n4219), .A2(n1212), .ZN(n6156) );
  INV_X2 U69 ( .A(n5732), .ZN(n5737) );
  INV_X2 U72 ( .A(n1691), .ZN(n771) );
  OAI22_X1 U76 ( .A1(n1129), .A2(n4100), .B1(n4108), .B2(n4101), .ZN(n1128) );
  NOR2_X2 U77 ( .A1(n3732), .A2(n5723), .ZN(n1692) );
  NOR2_X2 U79 ( .A1(n3317), .A2(n3361), .ZN(n5723) );
  INV_X4 U87 ( .A(n4199), .ZN(n6332) );
  NAND2_X1 U89 ( .A1(n4001), .A2(n1865), .ZN(n3810) );
  OR2_X2 U91 ( .A1(n1120), .A2(n2438), .ZN(n1452) );
  NAND2_X1 U100 ( .A1(n1120), .A2(n2438), .ZN(n1450) );
  NAND2_X2 U101 ( .A1(n5802), .A2(n5800), .ZN(n5801) );
  AND2_X2 U104 ( .A1(n2887), .A2(a[23]), .ZN(n6040) );
  XNOR2_X2 U114 ( .A(a[15]), .B(b[21]), .ZN(n5196) );
  XNOR2_X2 U116 ( .A(a[15]), .B(b[19]), .ZN(n5078) );
  XNOR2_X2 U118 ( .A(a[15]), .B(b[3]), .ZN(n3925) );
  XNOR2_X2 U119 ( .A(a[15]), .B(b[6]), .ZN(n4359) );
  NAND2_X2 U120 ( .A1(a[15]), .A2(n311), .ZN(n312) );
  XNOR2_X2 U125 ( .A(a[15]), .B(b[12]), .ZN(n4704) );
  XNOR2_X2 U133 ( .A(a[15]), .B(b[9]), .ZN(n4500) );
  NOR2_X2 U134 ( .A1(n501), .A2(a[15]), .ZN(n3394) );
  NAND2_X1 U143 ( .A1(n2384), .A2(n1844), .ZN(n1073) );
  NAND2_X2 U144 ( .A1(a[21]), .A2(n6515), .ZN(n3597) );
  NAND2_X1 U153 ( .A1(a[21]), .A2(n5360), .ZN(n3198) );
  NAND2_X1 U158 ( .A1(n981), .A2(a[21]), .ZN(n4992) );
  INV_X2 U165 ( .A(n4769), .ZN(n6658) );
  INV_X2 U166 ( .A(n4916), .ZN(n574) );
  NAND2_X2 U167 ( .A1(n5105), .A2(a[3]), .ZN(n4588) );
  INV_X2 U172 ( .A(n1239), .ZN(n653) );
  NAND2_X1 U188 ( .A1(n1239), .A2(n2824), .ZN(n655) );
  NOR2_X1 U193 ( .A1(n3639), .A2(a[11]), .ZN(n5100) );
  NAND2_X4 U200 ( .A1(n5718), .A2(n5717), .ZN(n2294) );
  AND2_X2 U204 ( .A1(n4358), .A2(n4357), .ZN(n6455) );
  NOR2_X2 U207 ( .A1(n1455), .A2(n3968), .ZN(n3345) );
  NOR2_X2 U210 ( .A1(n1455), .A2(n5002), .ZN(n1045) );
  NAND2_X1 U212 ( .A1(n3452), .A2(n3153), .ZN(n325) );
  NAND2_X4 U218 ( .A1(n6289), .A2(n6288), .ZN(n1089) );
  INV_X2 U219 ( .A(n3654), .ZN(n3937) );
  INV_X2 U220 ( .A(n5239), .ZN(n3231) );
  NAND2_X1 U221 ( .A1(n4910), .A2(n3608), .ZN(n210) );
  INV_X1 U227 ( .A(n2459), .ZN(n2458) );
  NAND2_X4 U231 ( .A1(n6284), .A2(n2546), .ZN(n1852) );
  INV_X4 U234 ( .A(n2767), .ZN(n2864) );
  NOR3_X2 U238 ( .A1(n5925), .A2(n2767), .A3(n5923), .ZN(n6111) );
  OAI21_X1 U242 ( .B1(n2765), .B2(n1850), .A(n4917), .ZN(n1952) );
  INV_X4 U243 ( .A(n6132), .ZN(n924) );
  NAND2_X4 U245 ( .A1(n3146), .A2(n1053), .ZN(n1360) );
  INV_X1 U260 ( .A(n2126), .ZN(n2091) );
  NAND2_X4 U262 ( .A1(n5108), .A2(n5107), .ZN(n5164) );
  NAND2_X4 U263 ( .A1(n3586), .A2(n5105), .ZN(n5108) );
  NAND2_X4 U265 ( .A1(n6026), .A2(n3540), .ZN(n4324) );
  NAND2_X1 U266 ( .A1(n146), .A2(n3073), .ZN(n1375) );
  NAND2_X1 U277 ( .A1(n2769), .A2(n3073), .ZN(n2693) );
  NAND2_X1 U279 ( .A1(n2773), .A2(n4719), .ZN(n779) );
  INV_X2 U288 ( .A(n3347), .ZN(n2368) );
  NOR2_X4 U291 ( .A1(n2282), .A2(n2281), .ZN(n4650) );
  NOR2_X4 U292 ( .A1(n6380), .A2(n2279), .ZN(n4651) );
  NAND2_X1 U293 ( .A1(n291), .A2(n2160), .ZN(n6270) );
  NAND2_X2 U295 ( .A1(n4092), .A2(a[5]), .ZN(n6456) );
  NAND2_X2 U303 ( .A1(n4092), .A2(a[5]), .ZN(n6457) );
  NAND2_X2 U309 ( .A1(n4933), .A2(n75), .ZN(n460) );
  NAND2_X1 U311 ( .A1(n4035), .A2(n4036), .ZN(n3594) );
  NAND2_X4 U316 ( .A1(n3542), .A2(n2225), .ZN(n3910) );
  NOR2_X1 U321 ( .A1(n1012), .A2(b[3]), .ZN(n6383) );
  OR2_X1 U322 ( .A1(n4543), .A2(b[17]), .ZN(n20) );
  NAND2_X2 U344 ( .A1(n4399), .A2(n585), .ZN(n4512) );
  NAND2_X2 U355 ( .A1(n1847), .A2(n984), .ZN(n4397) );
  INV_X2 U357 ( .A(n4972), .ZN(n3428) );
  NAND2_X2 U358 ( .A1(n1288), .A2(n6094), .ZN(n2894) );
  INV_X2 U359 ( .A(n1288), .ZN(n2892) );
  INV_X4 U362 ( .A(n6492), .ZN(n3427) );
  INV_X2 U367 ( .A(n5876), .ZN(n6509) );
  INV_X2 U370 ( .A(n5627), .ZN(n5626) );
  NAND2_X2 U371 ( .A1(n6453), .A2(n5813), .ZN(n5790) );
  INV_X2 U390 ( .A(n1666), .ZN(n191) );
  AND2_X2 U395 ( .A1(n3375), .A2(n5040), .ZN(n6461) );
  INV_X2 U396 ( .A(n3287), .ZN(n3286) );
  NAND2_X2 U400 ( .A1(n2552), .A2(n2551), .ZN(n4306) );
  NAND2_X2 U406 ( .A1(n904), .A2(n905), .ZN(n6440) );
  INV_X2 U414 ( .A(n6649), .ZN(n6449) );
  OR2_X2 U417 ( .A1(n6053), .A2(n6054), .ZN(n6469) );
  INV_X4 U428 ( .A(n4918), .ZN(n5039) );
  INV_X2 U433 ( .A(n2418), .ZN(n1642) );
  INV_X2 U434 ( .A(n2348), .ZN(n124) );
  NAND2_X2 U440 ( .A1(n2350), .A2(n2351), .ZN(n2349) );
  INV_X2 U441 ( .A(n4667), .ZN(n1030) );
  INV_X2 U450 ( .A(n1105), .ZN(n4196) );
  NAND2_X2 U466 ( .A1(n1463), .A2(n1462), .ZN(n3103) );
  INV_X2 U467 ( .A(n2258), .ZN(n6597) );
  NAND2_X2 U478 ( .A1(n3036), .A2(n3035), .ZN(n3040) );
  INV_X4 U488 ( .A(n2484), .ZN(n3510) );
  BUF_X2 U491 ( .A(n782), .Z(n185) );
  NAND2_X2 U495 ( .A1(n3736), .A2(n2925), .ZN(n2919) );
  OR2_X2 U505 ( .A1(n5295), .A2(n5294), .ZN(n6507) );
  NOR2_X2 U506 ( .A1(n6286), .A2(n6285), .ZN(n2216) );
  INV_X2 U507 ( .A(n4248), .ZN(n287) );
  INV_X2 U520 ( .A(n2616), .ZN(n2614) );
  NAND2_X2 U532 ( .A1(n3137), .A2(b[12]), .ZN(n238) );
  NAND2_X2 U545 ( .A1(n3692), .A2(n3691), .ZN(n3690) );
  INV_X4 U548 ( .A(n6566), .ZN(n3137) );
  INV_X8 U549 ( .A(n5197), .ZN(n6459) );
  INV_X4 U568 ( .A(n6479), .ZN(n938) );
  NAND2_X2 U570 ( .A1(n3793), .A2(a[13]), .ZN(n3791) );
  XOR2_X2 U571 ( .A(a[19]), .B(b[2]), .Z(n4428) );
  XOR2_X2 U573 ( .A(a[19]), .B(b[3]), .Z(n4349) );
  NOR2_X2 U574 ( .A1(a[9]), .A2(a[10]), .ZN(n6616) );
  NAND2_X2 U575 ( .A1(b[0]), .A2(a[1]), .ZN(n5642) );
  AND2_X2 U586 ( .A1(b[0]), .A2(a[0]), .ZN(\d[0] ) );
  INV_X4 U587 ( .A(n4924), .ZN(n6460) );
  XOR2_X2 U591 ( .A(a[3]), .B(b[5]), .Z(n1474) );
  INV_X4 U632 ( .A(b[13]), .ZN(n184) );
  XOR2_X2 U635 ( .A(a[13]), .B(b[2]), .Z(n3777) );
  XOR2_X2 U637 ( .A(a[3]), .B(b[15]), .Z(n3920) );
  XNOR2_X1 U638 ( .A(a[17]), .B(b[12]), .ZN(n4828) );
  NAND2_X1 U650 ( .A1(n699), .A2(n5529), .ZN(n2591) );
  NAND2_X1 U656 ( .A1(n4821), .A2(n3131), .ZN(n4537) );
  XNOR2_X1 U660 ( .A(b[10]), .B(a[19]), .ZN(n4825) );
  NAND3_X1 U661 ( .A1(n4835), .A2(n1062), .A3(n4724), .ZN(n4680) );
  INV_X2 U674 ( .A(n4678), .ZN(n4658) );
  INV_X1 U679 ( .A(n6605), .ZN(n4797) );
  NAND2_X1 U681 ( .A1(n4532), .A2(n4998), .ZN(n4533) );
  NOR2_X1 U685 ( .A1(n699), .A2(b[16]), .ZN(n1442) );
  NAND2_X1 U686 ( .A1(n1760), .A2(b[11]), .ZN(n4991) );
  NOR2_X1 U690 ( .A1(n5077), .A2(n5293), .ZN(n4787) );
  NAND2_X1 U705 ( .A1(n4835), .A2(n1062), .ZN(n4744) );
  INV_X2 U709 ( .A(n5015), .ZN(n5018) );
  XOR2_X1 U711 ( .A(b[18]), .B(a[3]), .Z(n2730) );
  NOR2_X2 U739 ( .A1(n5077), .A2(n3342), .ZN(n4501) );
  NAND2_X1 U742 ( .A1(n3431), .A2(n5360), .ZN(n3330) );
  INV_X1 U744 ( .A(n4926), .ZN(n301) );
  NAND2_X2 U745 ( .A1(n501), .A2(a[13]), .ZN(n504) );
  NAND2_X2 U751 ( .A1(n564), .A2(n2732), .ZN(n6620) );
  AOI22_X1 U757 ( .A1(n4705), .A2(b[6]), .B1(n1207), .B2(n1324), .ZN(n3921) );
  INV_X2 U758 ( .A(n2990), .ZN(n2897) );
  INV_X1 U759 ( .A(n2076), .ZN(n5111) );
  NAND2_X1 U760 ( .A1(n5109), .A2(n3540), .ZN(n3163) );
  NOR2_X1 U770 ( .A1(n4216), .A2(n4942), .ZN(n6234) );
  NAND2_X2 U787 ( .A1(n6304), .A2(n4330), .ZN(n6213) );
  NAND2_X1 U789 ( .A1(n5167), .A2(n5166), .ZN(n1205) );
  OAI21_X1 U793 ( .B1(n6203), .B2(n2249), .A(n2248), .ZN(n2247) );
  AOI21_X1 U802 ( .B1(n2844), .B2(n3747), .A(n3965), .ZN(n6488) );
  NAND2_X1 U806 ( .A1(n4913), .A2(n565), .ZN(n1382) );
  NOR2_X1 U807 ( .A1(n4284), .A2(n4283), .ZN(n4286) );
  INV_X2 U814 ( .A(n1003), .ZN(n6193) );
  NAND2_X2 U816 ( .A1(n1453), .A2(n1452), .ZN(n4294) );
  NAND2_X1 U818 ( .A1(n4648), .A2(n4649), .ZN(n1098) );
  INV_X2 U826 ( .A(n4085), .ZN(n3701) );
  INV_X2 U828 ( .A(n6086), .ZN(n6680) );
  NAND2_X1 U835 ( .A1(n4716), .A2(n4712), .ZN(n4714) );
  AND2_X2 U854 ( .A1(b[7]), .A2(b[6]), .ZN(n6462) );
  INV_X2 U860 ( .A(n4566), .ZN(n4565) );
  OR2_X2 U861 ( .A1(n2844), .A2(n3747), .ZN(n6463) );
  AND2_X2 U864 ( .A1(n6522), .A2(n2948), .ZN(n6464) );
  OR2_X2 U868 ( .A1(n2771), .A2(n1849), .ZN(n6465) );
  XOR2_X2 U873 ( .A(a[21]), .B(b[13]), .Z(n6466) );
  INV_X2 U874 ( .A(n1759), .ZN(n822) );
  AND2_X1 U875 ( .A1(b[7]), .A2(a[23]), .ZN(n6467) );
  INV_X1 U878 ( .A(n4906), .ZN(n3641) );
  OR2_X2 U882 ( .A1(n1682), .A2(n2447), .ZN(n6468) );
  INV_X2 U883 ( .A(n2141), .ZN(n6578) );
  NAND3_X2 U884 ( .A1(n2276), .A2(n3832), .A3(n3831), .ZN(n2141) );
  NAND2_X2 U900 ( .A1(n2427), .A2(n4282), .ZN(n2285) );
  NAND3_X2 U902 ( .A1(n2429), .A2(n2138), .A3(n2133), .ZN(n2427) );
  NAND2_X2 U903 ( .A1(n2646), .A2(n6470), .ZN(n4438) );
  NAND2_X1 U904 ( .A1(n1710), .A2(n4429), .ZN(n6470) );
  NAND2_X2 U905 ( .A1(n5395), .A2(n1547), .ZN(n5885) );
  NAND2_X2 U915 ( .A1(n5328), .A2(n5327), .ZN(n1547) );
  OAI22_X2 U927 ( .A1(n4746), .A2(b[3]), .B1(n3539), .B2(n4694), .ZN(n3833) );
  NAND3_X2 U933 ( .A1(n6617), .A2(n4507), .A3(n6558), .ZN(n1364) );
  OAI21_X2 U937 ( .B1(n4395), .B2(n4396), .A(n3327), .ZN(n6617) );
  OAI21_X1 U949 ( .B1(n6471), .B2(n3322), .A(n3967), .ZN(n6482) );
  INV_X2 U968 ( .A(n6472), .ZN(n6471) );
  NAND2_X2 U976 ( .A1(n2987), .A2(n2373), .ZN(n6472) );
  NAND2_X2 U982 ( .A1(n6473), .A2(n6581), .ZN(n5869) );
  INV_X2 U984 ( .A(n2067), .ZN(n6473) );
  NAND2_X2 U985 ( .A1(n1342), .A2(n1341), .ZN(n2067) );
  NOR2_X1 U990 ( .A1(n806), .A2(n5951), .ZN(n3505) );
  NAND3_X2 U991 ( .A1(n1384), .A2(a[13]), .A3(a[14]), .ZN(n806) );
  NOR2_X2 U993 ( .A1(n4438), .A2(n4449), .ZN(n4441) );
  NOR2_X2 U994 ( .A1(n2579), .A2(n5321), .ZN(n5768) );
  NAND2_X2 U1002 ( .A1(n1429), .A2(n1430), .ZN(n2579) );
  NAND3_X2 U1008 ( .A1(n6475), .A2(n3709), .A3(n6474), .ZN(n2222) );
  INV_X2 U1010 ( .A(n4367), .ZN(n6474) );
  INV_X2 U1011 ( .A(n4368), .ZN(n6475) );
  NAND2_X4 U1040 ( .A1(n6477), .A2(n6476), .ZN(n3604) );
  OAI21_X2 U1042 ( .B1(n3332), .B2(n2041), .A(n1710), .ZN(n6476) );
  NAND3_X2 U1047 ( .A1(n6169), .A2(n6168), .A3(n3255), .ZN(n6477) );
  NOR2_X4 U1054 ( .A1(n2708), .A2(n4636), .ZN(n6496) );
  NOR2_X4 U1057 ( .A1(n6496), .A2(n4480), .ZN(n1866) );
  NAND2_X2 U1065 ( .A1(n1843), .A2(n1842), .ZN(n6366) );
  NAND2_X2 U1071 ( .A1(n170), .A2(n6478), .ZN(n3232) );
  NAND3_X2 U1081 ( .A1(n2184), .A2(n4465), .A3(n4463), .ZN(n6478) );
  NAND2_X2 U1082 ( .A1(n4408), .A2(n4366), .ZN(n3709) );
  NOR2_X4 U1084 ( .A1(a[16]), .A2(a[15]), .ZN(n6479) );
  AOI22_X2 U1086 ( .A1(n1287), .A2(n4017), .B1(n2994), .B2(n3048), .ZN(n3070)
         );
  INV_X4 U1093 ( .A(n6480), .ZN(n798) );
  NOR2_X2 U1108 ( .A1(n1566), .A2(n4466), .ZN(n6480) );
  INV_X2 U1109 ( .A(n3947), .ZN(n3946) );
  XNOR2_X2 U1110 ( .A(n3944), .B(n3945), .ZN(n3947) );
  XNOR2_X2 U1117 ( .A(n3213), .B(n2387), .ZN(n2016) );
  NAND2_X2 U1121 ( .A1(n4009), .A2(n1257), .ZN(n3213) );
  NAND2_X2 U1125 ( .A1(n4422), .A2(n4544), .ZN(n4426) );
  INV_X4 U1139 ( .A(a[17]), .ZN(n4422) );
  NAND2_X2 U1149 ( .A1(n3260), .A2(n4652), .ZN(n3014) );
  NOR3_X2 U1150 ( .A1(n3761), .A2(n963), .A3(n4615), .ZN(n3260) );
  NAND3_X1 U1154 ( .A1(n6654), .A2(a[13]), .A3(n4614), .ZN(n6656) );
  NAND3_X2 U1161 ( .A1(n787), .A2(n4488), .A3(n1027), .ZN(n2119) );
  NAND2_X2 U1166 ( .A1(n5328), .A2(n5327), .ZN(n533) );
  NAND3_X2 U1176 ( .A1(n2007), .A2(n2903), .A3(n5323), .ZN(n5328) );
  INV_X4 U1179 ( .A(n4445), .ZN(n578) );
  NAND2_X2 U1182 ( .A1(n6481), .A2(n2220), .ZN(n1568) );
  NAND2_X2 U1183 ( .A1(n2222), .A2(n2221), .ZN(n6481) );
  AOI21_X2 U1185 ( .B1(n3097), .B2(n4636), .A(n2708), .ZN(n3448) );
  AOI22_X2 U1187 ( .A1(n6561), .A2(n5793), .B1(n452), .B2(n2374), .ZN(n1690)
         );
  NAND2_X2 U1200 ( .A1(n6482), .A2(n3122), .ZN(n4008) );
  NAND2_X2 U1208 ( .A1(n63), .A2(n4039), .ZN(n1893) );
  INV_X4 U1209 ( .A(n6483), .ZN(n250) );
  NOR2_X2 U1223 ( .A1(n2993), .A2(n3495), .ZN(n6483) );
  NAND3_X2 U1224 ( .A1(n2878), .A2(n6133), .A3(n3157), .ZN(n6136) );
  NAND2_X2 U1226 ( .A1(n3204), .A2(n1441), .ZN(n4782) );
  NOR2_X2 U1238 ( .A1(n3069), .A2(n3070), .ZN(n3043) );
  NAND2_X2 U1241 ( .A1(n3046), .A2(n3044), .ZN(n3069) );
  NAND3_X2 U1248 ( .A1(n5618), .A2(n5619), .A3(n152), .ZN(\d[40] ) );
  NAND2_X1 U1255 ( .A1(n1902), .A2(n2728), .ZN(n2807) );
  NAND2_X2 U1264 ( .A1(n1922), .A2(n3812), .ZN(n3987) );
  NAND2_X2 U1275 ( .A1(n6626), .A2(n6625), .ZN(n1922) );
  NAND3_X2 U1279 ( .A1(n5874), .A2(n5615), .A3(n5616), .ZN(n5618) );
  NAND2_X2 U1285 ( .A1(n6484), .A2(n6281), .ZN(n3219) );
  NAND2_X2 U1288 ( .A1(n355), .A2(n354), .ZN(n6484) );
  NAND3_X2 U1295 ( .A1(n4664), .A2(n6486), .A3(n6485), .ZN(n4719) );
  NAND2_X2 U1319 ( .A1(n5106), .A2(b[14]), .ZN(n6485) );
  INV_X2 U1327 ( .A(n6533), .ZN(n6486) );
  NAND3_X2 U1328 ( .A1(n5922), .A2(n5094), .A3(n6350), .ZN(n5096) );
  NOR2_X4 U1331 ( .A1(n5377), .A2(n5622), .ZN(n5922) );
  NAND3_X2 U1332 ( .A1(n2222), .A2(n2221), .A3(n4444), .ZN(n1567) );
  NAND2_X2 U1357 ( .A1(n3067), .A2(n4368), .ZN(n2221) );
  NAND2_X2 U1376 ( .A1(n5328), .A2(n5327), .ZN(n2908) );
  INV_X2 U1379 ( .A(n1662), .ZN(n300) );
  NAND2_X2 U1380 ( .A1(n167), .A2(n4927), .ZN(n1662) );
  INV_X2 U1388 ( .A(n3240), .ZN(n2890) );
  NAND2_X2 U1391 ( .A1(n6311), .A2(n456), .ZN(n3240) );
  NAND2_X2 U1394 ( .A1(n6379), .A2(n1319), .ZN(n908) );
  NAND3_X2 U1398 ( .A1(n1289), .A2(n3276), .A3(n3981), .ZN(n1319) );
  NOR2_X2 U1401 ( .A1(n1799), .A2(n2593), .ZN(n1798) );
  NAND2_X2 U1402 ( .A1(n1371), .A2(n6438), .ZN(n1799) );
  NAND2_X2 U1403 ( .A1(n6487), .A2(n6463), .ZN(n4044) );
  INV_X2 U1413 ( .A(n6488), .ZN(n6487) );
  NAND2_X2 U1418 ( .A1(n6587), .A2(n629), .ZN(n3089) );
  NAND2_X2 U1423 ( .A1(n303), .A2(n302), .ZN(n6587) );
  NAND2_X2 U1425 ( .A1(n131), .A2(n6489), .ZN(n3900) );
  NAND3_X1 U1431 ( .A1(n3185), .A2(n3186), .A3(n3910), .ZN(n6489) );
  NAND2_X2 U1433 ( .A1(n6620), .A2(n3744), .ZN(n6640) );
  NAND2_X2 U1437 ( .A1(n1932), .A2(n1933), .ZN(n3744) );
  NOR2_X2 U1438 ( .A1(n6490), .A2(n2263), .ZN(n131) );
  NOR2_X2 U1462 ( .A1(n3185), .A2(n3910), .ZN(n6490) );
  NAND2_X4 U1484 ( .A1(n2238), .A2(n1319), .ZN(n5735) );
  INV_X4 U1498 ( .A(n4010), .ZN(n6654) );
  INV_X8 U1517 ( .A(n6654), .ZN(n817) );
  NAND2_X2 U1552 ( .A1(n1078), .A2(n1077), .ZN(n528) );
  NAND2_X2 U1561 ( .A1(n6442), .A2(n2902), .ZN(n1078) );
  BUF_X4 U1579 ( .A(n5804), .Z(n6491) );
  NAND2_X2 U1601 ( .A1(n5395), .A2(n1547), .ZN(n6525) );
  NAND2_X2 U1606 ( .A1(n3670), .A2(n5863), .ZN(n6010) );
  NAND2_X2 U1609 ( .A1(n5098), .A2(n5097), .ZN(n5863) );
  NAND2_X4 U1612 ( .A1(n6010), .A2(n5998), .ZN(n256) );
  NAND2_X2 U1615 ( .A1(n3606), .A2(n3605), .ZN(n3754) );
  NAND2_X2 U1621 ( .A1(n6457), .A2(n5471), .ZN(n3605) );
  NAND2_X2 U1632 ( .A1(n5735), .A2(n5733), .ZN(n3274) );
  INV_X2 U1634 ( .A(n3745), .ZN(n6639) );
  INV_X2 U1635 ( .A(n5842), .ZN(n6492) );
  AOI21_X2 U1646 ( .B1(n6493), .B2(n1927), .A(n2307), .ZN(n3975) );
  INV_X2 U1652 ( .A(n6494), .ZN(n6493) );
  NOR2_X2 U1665 ( .A1(n6155), .A2(b[12]), .ZN(n6494) );
  NAND2_X4 U1666 ( .A1(n533), .A2(n5596), .ZN(n1902) );
  INV_X2 U1671 ( .A(n2977), .ZN(n925) );
  NAND2_X2 U1679 ( .A1(n5329), .A2(n256), .ZN(n2977) );
  NAND2_X2 U1680 ( .A1(n3900), .A2(n3901), .ZN(n3902) );
  NAND2_X2 U1682 ( .A1(n6672), .A2(n6620), .ZN(n3186) );
  INV_X4 U1683 ( .A(a[1]), .ZN(n6628) );
  NAND3_X1 U1684 ( .A1(n3123), .A2(n4044), .A3(n320), .ZN(n3122) );
  BUF_X4 U1687 ( .A(n4467), .Z(n6495) );
  NAND2_X2 U1688 ( .A1(n2913), .A2(n3201), .ZN(n1262) );
  OAI21_X2 U1703 ( .B1(n4521), .B2(n458), .A(n3571), .ZN(n3201) );
  OAI21_X2 U1709 ( .B1(n1298), .B2(n2310), .A(n3910), .ZN(n1295) );
  NAND2_X2 U1735 ( .A1(n3662), .A2(n3744), .ZN(n1298) );
  NOR2_X2 U1737 ( .A1(n337), .A2(n4070), .ZN(n4074) );
  NAND2_X2 U1744 ( .A1(n6497), .A2(n3095), .ZN(n2652) );
  NAND2_X2 U1745 ( .A1(n3500), .A2(n646), .ZN(n6497) );
  NAND2_X2 U1751 ( .A1(n2118), .A2(n6149), .ZN(n4582) );
  XNOR2_X2 U1761 ( .A(n6498), .B(n2722), .ZN(n4475) );
  AOI22_X2 U1762 ( .A1(n2224), .A2(n2542), .B1(n6191), .B2(n2543), .ZN(n6498)
         );
  NOR2_X2 U1769 ( .A1(n7), .A2(n4636), .ZN(n2034) );
  NAND2_X2 U1770 ( .A1(n6499), .A2(n380), .ZN(n4388) );
  NAND2_X2 U1771 ( .A1(n378), .A2(n379), .ZN(n6499) );
  INV_X2 U1778 ( .A(n6500), .ZN(n3049) );
  NAND2_X2 U1793 ( .A1(n3148), .A2(n1104), .ZN(n6500) );
  NAND3_X2 U1797 ( .A1(n6174), .A2(n4325), .A3(n776), .ZN(n4486) );
  NAND2_X2 U1798 ( .A1(n6592), .A2(n291), .ZN(n4325) );
  NAND2_X2 U1799 ( .A1(n6501), .A2(n579), .ZN(n1566) );
  NAND2_X2 U1811 ( .A1(n578), .A2(n577), .ZN(n6501) );
  NAND2_X2 U1813 ( .A1(n6503), .A2(n6502), .ZN(n4341) );
  NAND2_X2 U1823 ( .A1(n512), .A2(n981), .ZN(n6502) );
  NAND2_X2 U1825 ( .A1(n1354), .A2(b[11]), .ZN(n6503) );
  INV_X4 U1833 ( .A(n4306), .ZN(n6504) );
  NAND2_X2 U1846 ( .A1(n4219), .A2(n6221), .ZN(n4220) );
  NAND2_X1 U1847 ( .A1(n6552), .A2(n901), .ZN(n6505) );
  AOI21_X1 U1848 ( .B1(n3996), .B2(n1552), .A(n921), .ZN(n1551) );
  NAND2_X1 U1850 ( .A1(n3219), .A2(n3641), .ZN(n879) );
  NAND2_X1 U1852 ( .A1(n2032), .A2(n2954), .ZN(n5071) );
  NAND2_X2 U1854 ( .A1(n1543), .A2(n1544), .ZN(n6506) );
  NAND2_X2 U1870 ( .A1(n1543), .A2(n1544), .ZN(n3134) );
  NAND3_X1 U1892 ( .A1(n4982), .A2(n4977), .A3(n2976), .ZN(n4983) );
  NAND2_X1 U1900 ( .A1(n2960), .A2(n4759), .ZN(n2959) );
  NOR2_X1 U1902 ( .A1(n3573), .A2(n950), .ZN(n1921) );
  NAND2_X1 U1904 ( .A1(n2834), .A2(n1215), .ZN(n2192) );
  INV_X2 U1916 ( .A(n3608), .ZN(n788) );
  NAND2_X1 U1920 ( .A1(n1560), .A2(n1711), .ZN(n894) );
  NAND2_X1 U1923 ( .A1(n5304), .A2(n5305), .ZN(n5353) );
  NAND2_X1 U1937 ( .A1(n1730), .A2(n6507), .ZN(n6508) );
  NAND2_X2 U1938 ( .A1(n1730), .A2(n6507), .ZN(n5369) );
  INV_X2 U1952 ( .A(n6071), .ZN(n5876) );
  INV_X1 U1953 ( .A(n5564), .ZN(n1100) );
  AOI22_X1 U1967 ( .A1(n2224), .A2(n2542), .B1(n6191), .B2(n2543), .ZN(n6510)
         );
  INV_X2 U1970 ( .A(n1049), .ZN(n2542) );
  INV_X4 U1975 ( .A(n5459), .ZN(n385) );
  NAND2_X2 U1977 ( .A1(n303), .A2(n302), .ZN(n4960) );
  NAND3_X2 U1994 ( .A1(n1480), .A2(n209), .A3(n1478), .ZN(n6511) );
  NAND2_X2 U1995 ( .A1(n2500), .A2(n2849), .ZN(n6512) );
  INV_X4 U1999 ( .A(n2503), .ZN(n6513) );
  NAND2_X1 U2001 ( .A1(n4504), .A2(b[3]), .ZN(n6550) );
  NOR2_X1 U2003 ( .A1(n4504), .A2(n4598), .ZN(n6243) );
  INV_X1 U2004 ( .A(n1710), .ZN(n6168) );
  INV_X2 U2006 ( .A(n680), .ZN(n4716) );
  NAND2_X2 U2031 ( .A1(n825), .A2(n826), .ZN(n6514) );
  INV_X4 U2044 ( .A(n2478), .ZN(n825) );
  NAND2_X1 U2045 ( .A1(n4904), .A2(n4903), .ZN(n6281) );
  INV_X1 U2057 ( .A(n4903), .ZN(n4905) );
  MUX2_X2 U2067 ( .A(n5899), .B(n6035), .S(n6515), .Z(n5444) );
  NAND2_X2 U2104 ( .A1(n1285), .A2(n1284), .ZN(n6516) );
  NAND2_X2 U2107 ( .A1(n1285), .A2(n1284), .ZN(n2044) );
  NAND2_X4 U2110 ( .A1(a[16]), .A2(a[15]), .ZN(n6517) );
  NAND2_X4 U2135 ( .A1(a[16]), .A2(a[15]), .ZN(n6518) );
  NAND2_X2 U2139 ( .A1(n5195), .A2(n5194), .ZN(n5226) );
  NOR2_X4 U2148 ( .A1(n5932), .A2(n5871), .ZN(n5996) );
  NAND2_X1 U2154 ( .A1(n6155), .A2(n184), .ZN(n92) );
  NAND2_X1 U2157 ( .A1(n6155), .A2(n3538), .ZN(n6387) );
  NAND2_X1 U2160 ( .A1(n6155), .A2(n4942), .ZN(n6318) );
  NAND2_X1 U2168 ( .A1(n6155), .A2(n4598), .ZN(n198) );
  INV_X4 U2173 ( .A(n477), .ZN(n4711) );
  NAND2_X2 U2180 ( .A1(n5928), .A2(n6134), .ZN(n6519) );
  NAND2_X2 U2183 ( .A1(n372), .A2(n373), .ZN(n6520) );
  NAND3_X1 U2184 ( .A1(n2953), .A2(n3698), .A3(n5182), .ZN(n2206) );
  NAND2_X1 U2191 ( .A1(n1521), .A2(n1522), .ZN(n565) );
  NAND2_X1 U2203 ( .A1(n6256), .A2(n3629), .ZN(n6521) );
  NOR2_X1 U2204 ( .A1(n5729), .A2(n3396), .ZN(n6522) );
  INV_X8 U2206 ( .A(n2037), .ZN(n5477) );
  NAND2_X1 U2209 ( .A1(n2532), .A2(n3318), .ZN(n6523) );
  NAND2_X2 U2212 ( .A1(n2532), .A2(n3318), .ZN(n1945) );
  NAND2_X2 U2225 ( .A1(n6056), .A2(n5631), .ZN(n5632) );
  NAND2_X1 U2228 ( .A1(n1761), .A2(n184), .ZN(n183) );
  AOI22_X2 U2237 ( .A1(n558), .A2(b[5]), .B1(n3835), .B2(n4940), .ZN(n2533) );
  NAND2_X4 U2239 ( .A1(n1893), .A2(n1892), .ZN(n2987) );
  INV_X1 U2249 ( .A(n328), .ZN(n6524) );
  NOR2_X2 U2250 ( .A1(n4069), .A2(n4068), .ZN(n4464) );
  INV_X4 U2255 ( .A(n1265), .ZN(n1264) );
  NAND2_X1 U2263 ( .A1(n558), .A2(b[23]), .ZN(n5223) );
  NAND2_X1 U2266 ( .A1(n558), .A2(b[19]), .ZN(n5000) );
  NAND2_X1 U2277 ( .A1(n1891), .A2(n4038), .ZN(n335) );
  INV_X2 U2281 ( .A(n1891), .ZN(n333) );
  NOR2_X1 U2282 ( .A1(b[14]), .A2(n3011), .ZN(n6533) );
  NAND2_X1 U2284 ( .A1(n984), .A2(n5266), .ZN(n6427) );
  OAI21_X1 U2285 ( .B1(n4377), .B2(n4376), .A(n4375), .ZN(n711) );
  NAND2_X2 U2289 ( .A1(n1278), .A2(n3568), .ZN(n1200) );
  NOR3_X2 U2301 ( .A1(n5968), .A2(n5628), .A3(n5971), .ZN(n6526) );
  NOR3_X2 U2311 ( .A1(n5968), .A2(n5628), .A3(n5971), .ZN(n5929) );
  NAND2_X4 U2312 ( .A1(a[4]), .A2(a[3]), .ZN(n6527) );
  NAND2_X4 U2313 ( .A1(a[4]), .A2(a[3]), .ZN(n6528) );
  INV_X2 U2314 ( .A(n6528), .ZN(n3435) );
  AOI22_X2 U2316 ( .A1(n4489), .A2(n3576), .B1(n4408), .B2(n3765), .ZN(n6529)
         );
  AOI22_X1 U2317 ( .A1(n4489), .A2(n3576), .B1(n4408), .B2(n3765), .ZN(n3199)
         );
  XOR2_X1 U2318 ( .A(n6510), .B(n2722), .Z(n6530) );
  AND2_X4 U2319 ( .A1(n4386), .A2(n4385), .ZN(n2722) );
  INV_X4 U2325 ( .A(n6531), .ZN(n6536) );
  NOR2_X2 U2326 ( .A1(n2005), .A2(n2004), .ZN(n6531) );
  NAND2_X2 U2327 ( .A1(n6532), .A2(n1232), .ZN(n1959) );
  NAND2_X2 U2332 ( .A1(n2399), .A2(n1960), .ZN(n6532) );
  NAND2_X2 U2333 ( .A1(n3509), .A2(n3346), .ZN(n3082) );
  NAND2_X2 U2339 ( .A1(n1832), .A2(n6644), .ZN(n3346) );
  NAND3_X1 U2355 ( .A1(n5998), .A2(n5596), .A3(n533), .ZN(n5329) );
  AOI22_X2 U2360 ( .A1(n4722), .A2(n4718), .B1(n4721), .B2(n4663), .ZN(n4904)
         );
  NOR2_X4 U2386 ( .A1(n6534), .A2(n1790), .ZN(n4759) );
  AOI22_X2 U2389 ( .A1(n2656), .A2(n981), .B1(n5336), .B2(b[11]), .ZN(n6534)
         );
  NAND2_X4 U2395 ( .A1(n6536), .A2(n6535), .ZN(n5860) );
  NAND2_X2 U2406 ( .A1(n2005), .A2(n2004), .ZN(n6535) );
  NAND2_X2 U2409 ( .A1(n6537), .A2(n570), .ZN(n572) );
  INV_X2 U2412 ( .A(n1083), .ZN(n6537) );
  NAND2_X2 U2413 ( .A1(n576), .A2(n575), .ZN(n1083) );
  INV_X2 U2417 ( .A(n6538), .ZN(n2254) );
  NOR2_X2 U2421 ( .A1(n1761), .A2(b[8]), .ZN(n6538) );
  OAI22_X2 U2425 ( .A1(n2950), .A2(n4598), .B1(n5266), .B2(b[4]), .ZN(n2271)
         );
  NAND2_X2 U2432 ( .A1(n6539), .A2(n6279), .ZN(n1691) );
  INV_X2 U2433 ( .A(n6540), .ZN(n6539) );
  NAND3_X2 U2435 ( .A1(n1340), .A2(n2364), .A3(n2294), .ZN(n6540) );
  NAND2_X2 U2436 ( .A1(n6020), .A2(n6541), .ZN(n6635) );
  AOI22_X2 U2441 ( .A1(n6018), .A2(n6019), .B1(n6021), .B2(n2822), .ZN(n6541)
         );
  NAND3_X2 U2443 ( .A1(n1939), .A2(n1938), .A3(n6542), .ZN(n1466) );
  INV_X2 U2448 ( .A(n4684), .ZN(n6542) );
  NOR2_X2 U2456 ( .A1(n4682), .A2(n4683), .ZN(n4684) );
  OAI21_X2 U2476 ( .B1(n3268), .B2(n4672), .A(n2216), .ZN(n1939) );
  NAND2_X2 U2504 ( .A1(n6613), .A2(n5858), .ZN(n2933) );
  NOR2_X4 U2516 ( .A1(n5851), .A2(n5854), .ZN(n6613) );
  NAND3_X2 U2529 ( .A1(n2144), .A2(n6591), .A3(n3171), .ZN(n1581) );
  AOI21_X1 U2538 ( .B1(n6336), .B2(n5834), .A(n2006), .ZN(n289) );
  NAND2_X2 U2540 ( .A1(n1573), .A2(n1572), .ZN(n4628) );
  NAND2_X2 U2559 ( .A1(n85), .A2(n84), .ZN(n1573) );
  NAND2_X2 U2565 ( .A1(n3520), .A2(n5823), .ZN(n2006) );
  NAND2_X2 U2604 ( .A1(n3234), .A2(n3235), .ZN(n4576) );
  XNOR2_X2 U2612 ( .A(n1333), .B(n2792), .ZN(n3235) );
  NAND2_X2 U2618 ( .A1(n677), .A2(n676), .ZN(n6336) );
  NAND2_X2 U2668 ( .A1(n6543), .A2(n2754), .ZN(n5029) );
  NAND3_X2 U2669 ( .A1(n3312), .A2(n4925), .A3(n1888), .ZN(n6543) );
  NAND2_X2 U2671 ( .A1(n6545), .A2(n6544), .ZN(n4597) );
  NAND2_X2 U2683 ( .A1(n5077), .A2(b[10]), .ZN(n6544) );
  NAND2_X2 U2703 ( .A1(n5076), .A2(n4942), .ZN(n6545) );
  NOR2_X4 U2711 ( .A1(n5477), .A2(n4752), .ZN(n4605) );
  NAND2_X4 U2713 ( .A1(n2038), .A2(a[23]), .ZN(n2037) );
  NAND4_X1 U2721 ( .A1(n2804), .A2(n324), .A3(n1581), .A4(n1028), .ZN(n563) );
  NOR3_X2 U2743 ( .A1(n5845), .A2(n3427), .A3(n5841), .ZN(n5847) );
  NAND2_X2 U2748 ( .A1(n1999), .A2(n2729), .ZN(n2855) );
  NOR2_X4 U2750 ( .A1(n6547), .A2(n6546), .ZN(n1999) );
  INV_X4 U2774 ( .A(n6517), .ZN(n6546) );
  INV_X4 U2800 ( .A(n938), .ZN(n6547) );
  NAND2_X4 U2807 ( .A1(n2472), .A2(n6572), .ZN(n2825) );
  INV_X4 U2816 ( .A(n6669), .ZN(n6165) );
  NAND2_X2 U2824 ( .A1(n6548), .A2(n6334), .ZN(n5665) );
  NAND2_X2 U2826 ( .A1(n6332), .A2(n6333), .ZN(n6548) );
  NAND2_X4 U2838 ( .A1(n938), .A2(n6518), .ZN(n2854) );
  NAND2_X2 U2844 ( .A1(n3564), .A2(n6549), .ZN(n2519) );
  NAND3_X1 U2856 ( .A1(n4187), .A2(n2508), .A3(n4231), .ZN(n6549) );
  NAND2_X2 U2870 ( .A1(n6551), .A2(n6550), .ZN(n4089) );
  NAND2_X1 U2880 ( .A1(n3431), .A2(n3538), .ZN(n6551) );
  NAND2_X2 U2882 ( .A1(n6552), .A2(n901), .ZN(n4312) );
  NAND2_X2 U2912 ( .A1(n899), .A2(n4302), .ZN(n6552) );
  NAND2_X1 U2922 ( .A1(n3517), .A2(n5282), .ZN(n2664) );
  NAND2_X2 U2924 ( .A1(n2661), .A2(n2660), .ZN(n3517) );
  NAND2_X4 U2934 ( .A1(n873), .A2(n6553), .ZN(n876) );
  INV_X2 U2944 ( .A(n1685), .ZN(n6553) );
  XNOR2_X2 U2945 ( .A(n4102), .B(n4101), .ZN(n1685) );
  NAND2_X2 U2966 ( .A1(n368), .A2(n1148), .ZN(n2452) );
  NAND2_X2 U2973 ( .A1(n1524), .A2(n164), .ZN(n3385) );
  NAND2_X2 U2975 ( .A1(n2449), .A2(n6277), .ZN(n1666) );
  NAND2_X2 U2976 ( .A1(n6555), .A2(n6554), .ZN(n1176) );
  INV_X2 U3006 ( .A(n3984), .ZN(n6554) );
  INV_X2 U3013 ( .A(n1175), .ZN(n6555) );
  NAND2_X2 U3019 ( .A1(n5578), .A2(n5579), .ZN(n5609) );
  NAND2_X2 U3020 ( .A1(n228), .A2(n623), .ZN(n5578) );
  NOR2_X2 U3022 ( .A1(n6556), .A2(n5874), .ZN(n1339) );
  NAND3_X2 U3040 ( .A1(n6525), .A2(n5878), .A3(n5872), .ZN(n6556) );
  INV_X4 U3061 ( .A(n2401), .ZN(n3384) );
  NAND2_X2 U3062 ( .A1(n5115), .A2(n5116), .ZN(n2401) );
  NAND2_X2 U3065 ( .A1(n3294), .A2(n4836), .ZN(n4837) );
  NAND2_X2 U3070 ( .A1(n3295), .A2(n3296), .ZN(n3294) );
  AOI22_X2 U3096 ( .A1(n6439), .A2(b[2]), .B1(n998), .B2(n2249), .ZN(n1208) );
  INV_X4 U3097 ( .A(n3524), .ZN(n1640) );
  NAND2_X2 U3110 ( .A1(n4995), .A2(n184), .ZN(n3692) );
  INV_X2 U3118 ( .A(n6557), .ZN(n3377) );
  NAND2_X2 U3123 ( .A1(n2600), .A2(n2599), .ZN(n6557) );
  AOI22_X2 U3132 ( .A1(n5900), .A2(b[7]), .B1(n435), .B2(n3465), .ZN(n4890) );
  NAND2_X2 U3133 ( .A1(n3090), .A2(n3089), .ZN(n487) );
  OAI21_X2 U3139 ( .B1(n4960), .B2(n629), .A(n1831), .ZN(n3090) );
  AOI22_X2 U3147 ( .A1(n5454), .A2(b[13]), .B1(n314), .B2(n4614), .ZN(n3323)
         );
  NAND2_X4 U3153 ( .A1(n3506), .A2(n4422), .ZN(n5454) );
  NAND3_X2 U3171 ( .A1(n4371), .A2(n3306), .A3(n3307), .ZN(n4373) );
  BUF_X4 U3172 ( .A(n6528), .Z(n6558) );
  NAND2_X2 U3174 ( .A1(n6559), .A2(n5126), .ZN(n5208) );
  INV_X2 U3180 ( .A(n5129), .ZN(n6559) );
  NAND2_X2 U3181 ( .A1(n1631), .A2(n1630), .ZN(n5129) );
  NAND2_X2 U3199 ( .A1(n6560), .A2(n4354), .ZN(n1575) );
  AOI22_X2 U3210 ( .A1(n1127), .A2(n4346), .B1(n4347), .B2(n4348), .ZN(n6560)
         );
  NAND2_X2 U3215 ( .A1(n5122), .A2(n1804), .ZN(n1815) );
  OAI22_X2 U3216 ( .A1(n2363), .A2(n2362), .B1(n2361), .B2(n5084), .ZN(n5122)
         );
  NAND2_X2 U3229 ( .A1(n2900), .A2(n4638), .ZN(n6561) );
  NAND2_X4 U3237 ( .A1(n6563), .A2(n6562), .ZN(n2175) );
  INV_X4 U3238 ( .A(n2177), .ZN(n6562) );
  INV_X4 U3248 ( .A(n1278), .ZN(n6563) );
  NAND2_X2 U3255 ( .A1(n4347), .A2(n4348), .ZN(n201) );
  NAND3_X2 U3262 ( .A1(n6564), .A2(n2141), .A3(n4270), .ZN(n2136) );
  NAND2_X2 U3278 ( .A1(n2275), .A2(n2274), .ZN(n6564) );
  NAND2_X2 U3283 ( .A1(a[5]), .A2(n6528), .ZN(n4789) );
  NAND2_X2 U3287 ( .A1(n5162), .A2(n2422), .ZN(n5099) );
  NAND2_X2 U3296 ( .A1(n6461), .A2(n2425), .ZN(n5162) );
  NAND2_X2 U3302 ( .A1(n4791), .A2(n4119), .ZN(n4104) );
  NAND2_X1 U3303 ( .A1(n4979), .A2(n4976), .ZN(n57) );
  XNOR2_X2 U3304 ( .A(n6565), .B(n3493), .ZN(n4275) );
  NAND2_X2 U3305 ( .A1(n1825), .A2(n1826), .ZN(n6565) );
  OAI21_X2 U3350 ( .B1(n1183), .B2(n3074), .A(n5039), .ZN(n3375) );
  INV_X2 U3352 ( .A(n3581), .ZN(n6566) );
  NAND2_X1 U3353 ( .A1(n1587), .A2(n28), .ZN(n6386) );
  NOR2_X2 U3363 ( .A1(n6568), .A2(n6567), .ZN(n28) );
  NOR2_X2 U3365 ( .A1(n3598), .A2(n4830), .ZN(n6567) );
  NOR2_X2 U3366 ( .A1(n4832), .A2(n4831), .ZN(n6568) );
  NOR2_X2 U3381 ( .A1(n4446), .A2(n2648), .ZN(n1565) );
  NOR2_X2 U3382 ( .A1(n4343), .A2(n15), .ZN(n4446) );
  NAND3_X2 U3389 ( .A1(n1017), .A2(n1752), .A3(n1753), .ZN(n1595) );
  OAI22_X2 U3395 ( .A1(n4074), .A2(n4073), .B1(n4071), .B2(n4072), .ZN(n4076)
         );
  BUF_X4 U3398 ( .A(n4544), .Z(n6569) );
  BUF_X4 U3399 ( .A(n4624), .Z(n6570) );
  NAND2_X2 U3400 ( .A1(n2793), .A2(n2272), .ZN(n4563) );
  NOR2_X2 U3421 ( .A1(n2621), .A2(n451), .ZN(n6285) );
  NAND2_X2 U3422 ( .A1(n6668), .A2(n6571), .ZN(n2993) );
  NAND3_X2 U3425 ( .A1(n6404), .A2(n470), .A3(n2925), .ZN(n6571) );
  OAI22_X2 U3429 ( .A1(n2147), .A2(n5190), .B1(n4605), .B2(n2603), .ZN(n4568)
         );
  OAI22_X2 U3430 ( .A1(n760), .A2(n3342), .B1(n6326), .B2(b[8]), .ZN(n6572) );
  NAND2_X2 U3448 ( .A1(n6574), .A2(n6573), .ZN(n1519) );
  INV_X2 U3449 ( .A(n1795), .ZN(n6573) );
  NAND2_X2 U3465 ( .A1(n2572), .A2(n2571), .ZN(n6574) );
  AOI21_X2 U3466 ( .B1(n2712), .B2(n2806), .A(n511), .ZN(n2805) );
  NAND2_X2 U3467 ( .A1(n6576), .A2(n6575), .ZN(n2712) );
  INV_X2 U3476 ( .A(n4555), .ZN(n6575) );
  INV_X2 U3481 ( .A(n4554), .ZN(n6576) );
  OAI21_X2 U3482 ( .B1(n4150), .B2(n5660), .A(n4149), .ZN(n3511) );
  NAND2_X2 U3488 ( .A1(n5657), .A2(n5658), .ZN(n4149) );
  NOR3_X2 U3489 ( .A1(n4147), .A2(n4146), .A3(n5658), .ZN(n4150) );
  NAND2_X2 U3522 ( .A1(n6577), .A2(n6399), .ZN(n2051) );
  INV_X2 U3524 ( .A(n5082), .ZN(n6577) );
  NOR2_X2 U3525 ( .A1(n6664), .A2(n4993), .ZN(n5082) );
  INV_X2 U3528 ( .A(n4629), .ZN(n3338) );
  NAND2_X2 U3529 ( .A1(n2608), .A2(n1574), .ZN(n4629) );
  AOI22_X2 U3530 ( .A1(n4995), .A2(n6221), .B1(b[9]), .B2(n465), .ZN(n6414) );
  NOR2_X2 U3533 ( .A1(n2966), .A2(n971), .ZN(n6663) );
  XNOR2_X2 U3534 ( .A(n5251), .B(n5239), .ZN(n2966) );
  NAND3_X2 U3539 ( .A1(n6618), .A2(n3357), .A3(n4287), .ZN(n2551) );
  NAND2_X2 U3540 ( .A1(n1900), .A2(n1901), .ZN(n6618) );
  NAND2_X2 U3563 ( .A1(n6578), .A2(n2430), .ZN(n2134) );
  NAND2_X4 U3585 ( .A1(n6579), .A2(n448), .ZN(n4316) );
  NAND2_X2 U3588 ( .A1(n447), .A2(n446), .ZN(n6579) );
  AND2_X2 U3589 ( .A1(n57), .A2(n5094), .ZN(n996) );
  OAI21_X2 U3593 ( .B1(n1718), .B2(n2946), .A(n3335), .ZN(n2940) );
  NOR2_X2 U3609 ( .A1(n2947), .A2(n4584), .ZN(n2946) );
  NAND2_X2 U3613 ( .A1(n6613), .A2(n1015), .ZN(n5374) );
  NAND2_X2 U3636 ( .A1(n6580), .A2(n5626), .ZN(n3677) );
  NAND2_X2 U3637 ( .A1(n3390), .A2(n3678), .ZN(n6580) );
  NAND2_X2 U3677 ( .A1(n5384), .A2(n1099), .ZN(n1145) );
  NAND2_X4 U3686 ( .A1(n6611), .A2(n5808), .ZN(n5384) );
  AOI22_X2 U3693 ( .A1(b[10]), .A2(n5472), .B1(n5897), .B2(n4942), .ZN(n4919)
         );
  NAND2_X4 U3700 ( .A1(n586), .A2(a[21]), .ZN(n5897) );
  INV_X4 U3722 ( .A(n5885), .ZN(n5589) );
  NOR2_X2 U3757 ( .A1(n4246), .A2(n921), .ZN(n4248) );
  INV_X2 U3762 ( .A(n5567), .ZN(n6581) );
  NAND2_X2 U3787 ( .A1(n727), .A2(n728), .ZN(n5567) );
  NAND2_X2 U3793 ( .A1(n6582), .A2(n3481), .ZN(n1502) );
  INV_X2 U3796 ( .A(n6583), .ZN(n6582) );
  NOR2_X2 U3806 ( .A1(n4590), .A2(n3263), .ZN(n6583) );
  INV_X2 U3823 ( .A(n6584), .ZN(n987) );
  NOR2_X2 U3829 ( .A1(n4893), .A2(n1531), .ZN(n6584) );
  INV_X4 U3842 ( .A(n6650), .ZN(n956) );
  NAND3_X1 U3843 ( .A1(n2635), .A2(n3250), .A3(n1146), .ZN(n3248) );
  NAND2_X2 U3853 ( .A1(n1689), .A2(n4731), .ZN(n2635) );
  NAND2_X2 U3879 ( .A1(n6374), .A2(n6373), .ZN(n5660) );
  BUF_X4 U3900 ( .A(n5947), .Z(n6585) );
  NOR2_X2 U3910 ( .A1(n6586), .A2(n4108), .ZN(n4117) );
  INV_X8 U3917 ( .A(n451), .ZN(n3308) );
  INV_X4 U3923 ( .A(n3026), .ZN(n2024) );
  NAND2_X4 U3931 ( .A1(n4213), .A2(n4214), .ZN(n4244) );
  NAND2_X1 U3947 ( .A1(n2045), .A2(n938), .ZN(n6588) );
  INV_X4 U3963 ( .A(n2829), .ZN(n6589) );
  INV_X2 U3966 ( .A(n3833), .ZN(n2276) );
  INV_X4 U3972 ( .A(n3843), .ZN(n3844) );
  INV_X4 U3979 ( .A(n4303), .ZN(n899) );
  NAND2_X2 U3999 ( .A1(n2021), .A2(n1305), .ZN(n6590) );
  NOR2_X1 U4000 ( .A1(n4175), .A2(n1626), .ZN(n5670) );
  NAND2_X1 U4002 ( .A1(n3235), .A2(n3234), .ZN(n6591) );
  NAND2_X1 U4025 ( .A1(n564), .A2(n2732), .ZN(n3662) );
  INV_X2 U4027 ( .A(n2160), .ZN(n6592) );
  AND2_X4 U4031 ( .A1(n2524), .A2(b[0]), .ZN(n2042) );
  NAND2_X1 U4032 ( .A1(n490), .A2(n491), .ZN(n6593) );
  NAND2_X2 U4036 ( .A1(n2017), .A2(n2018), .ZN(n6594) );
  NAND2_X2 U4041 ( .A1(n6595), .A2(n1286), .ZN(n4059) );
  INV_X2 U4044 ( .A(n6594), .ZN(n6595) );
  NAND2_X2 U4054 ( .A1(n6211), .A2(b[14]), .ZN(n2018) );
  INV_X2 U4055 ( .A(n4059), .ZN(n4065) );
  NOR2_X4 U4074 ( .A1(n3642), .A2(n4611), .ZN(n4672) );
  NAND2_X2 U4079 ( .A1(n4672), .A2(n6358), .ZN(n3290) );
  BUF_X4 U4081 ( .A(n4633), .Z(n6402) );
  NAND2_X1 U4087 ( .A1(n1200), .A2(n1197), .ZN(n6596) );
  NAND2_X1 U4091 ( .A1(n2258), .A2(n2257), .ZN(n6599) );
  NAND2_X2 U4111 ( .A1(n6597), .A2(n6598), .ZN(n6600) );
  NAND2_X2 U4116 ( .A1(n6599), .A2(n6600), .ZN(n3650) );
  INV_X1 U4125 ( .A(n2257), .ZN(n6598) );
  INV_X1 U4130 ( .A(n3911), .ZN(n2257) );
  NAND2_X2 U4139 ( .A1(n6590), .A2(n4975), .ZN(n6601) );
  NAND3_X2 U4140 ( .A1(n4026), .A2(a[18]), .A3(a[17]), .ZN(n465) );
  NOR2_X2 U4141 ( .A1(a[18]), .A2(a[17]), .ZN(n610) );
  NAND2_X2 U4153 ( .A1(a[18]), .A2(b[1]), .ZN(n4423) );
  INV_X4 U4156 ( .A(a[18]), .ZN(n4027) );
  INV_X1 U4194 ( .A(n610), .ZN(n4030) );
  NAND2_X1 U4204 ( .A1(n5179), .A2(b[3]), .ZN(n2617) );
  NAND2_X1 U4224 ( .A1(n5523), .A2(n5522), .ZN(n5892) );
  NAND2_X1 U4248 ( .A1(n5466), .A2(b[16]), .ZN(n5145) );
  NAND2_X1 U4250 ( .A1(n5466), .A2(b[15]), .ZN(n3623) );
  NAND3_X2 U4254 ( .A1(n4026), .A2(a[18]), .A3(a[17]), .ZN(n5179) );
  INV_X4 U4262 ( .A(n2033), .ZN(n6602) );
  INV_X2 U4269 ( .A(n2033), .ZN(n5798) );
  NAND2_X4 U4279 ( .A1(n245), .A2(n6353), .ZN(n3130) );
  INV_X1 U4281 ( .A(n4646), .ZN(n6603) );
  INV_X2 U4297 ( .A(n6603), .ZN(n6604) );
  INV_X2 U4305 ( .A(n4557), .ZN(n4646) );
  INV_X8 U4308 ( .A(a[6]), .ZN(n6606) );
  NAND2_X2 U4309 ( .A1(n1138), .A2(n4228), .ZN(n3564) );
  NOR2_X4 U4327 ( .A1(n2486), .A2(n2487), .ZN(n4503) );
  NAND2_X1 U4328 ( .A1(n4293), .A2(n4294), .ZN(n696) );
  NAND2_X2 U4329 ( .A1(n807), .A2(n2149), .ZN(n6607) );
  NAND2_X4 U4342 ( .A1(n674), .A2(n675), .ZN(n677) );
  INV_X4 U4345 ( .A(n6329), .ZN(n1654) );
  INV_X2 U4348 ( .A(n4060), .ZN(n4063) );
  NAND2_X2 U4350 ( .A1(n3264), .A2(n4526), .ZN(n2479) );
  NAND2_X4 U4383 ( .A1(n6440), .A2(n906), .ZN(n5681) );
  INV_X2 U4385 ( .A(n3264), .ZN(n3063) );
  NAND2_X2 U4404 ( .A1(n3638), .A2(n4998), .ZN(n3637) );
  INV_X2 U4422 ( .A(n3627), .ZN(n515) );
  NAND2_X1 U4424 ( .A1(n1387), .A2(n3727), .ZN(n4718) );
  OAI21_X1 U4434 ( .B1(n2195), .B2(n3887), .A(n2437), .ZN(n1404) );
  INV_X4 U4436 ( .A(n3603), .ZN(n98) );
  NOR2_X4 U4437 ( .A1(n4766), .A2(n3383), .ZN(n3603) );
  MUX2_X2 U4444 ( .A(n512), .B(n606), .S(b[5]), .Z(n3816) );
  NAND2_X2 U4446 ( .A1(n2586), .A2(n2585), .ZN(n6608) );
  NAND2_X2 U4450 ( .A1(b[18]), .A2(n2244), .ZN(n3644) );
  NAND2_X2 U4452 ( .A1(n2126), .A2(n2125), .ZN(n6609) );
  NAND2_X2 U4453 ( .A1(n2125), .A2(n2126), .ZN(n3731) );
  INV_X2 U4455 ( .A(n3015), .ZN(n2125) );
  INV_X2 U4461 ( .A(n3831), .ZN(n2274) );
  INV_X4 U4462 ( .A(n4613), .ZN(n4562) );
  NAND2_X2 U4465 ( .A1(n4352), .A2(n4353), .ZN(n6610) );
  NAND2_X2 U4466 ( .A1(n4353), .A2(n4352), .ZN(n4403) );
  INV_X4 U4489 ( .A(n5842), .ZN(n6611) );
  INV_X2 U4495 ( .A(n5798), .ZN(n5781) );
  NAND2_X2 U4501 ( .A1(n1125), .A2(n1122), .ZN(n906) );
  INV_X2 U4502 ( .A(n1560), .ZN(n892) );
  XNOR2_X2 U4503 ( .A(n6612), .B(b[23]), .ZN(n4586) );
  INV_X8 U4504 ( .A(a[3]), .ZN(n6612) );
  NOR2_X4 U4518 ( .A1(a[11]), .A2(a[12]), .ZN(n6614) );
  OR2_X2 U4525 ( .A1(n502), .A2(a[12]), .ZN(n953) );
  INV_X8 U4539 ( .A(a[12]), .ZN(n187) );
  NAND2_X1 U4548 ( .A1(n3803), .A2(n397), .ZN(n3804) );
  NOR2_X4 U4555 ( .A1(a[9]), .A2(a[10]), .ZN(n6615) );
  INV_X2 U4557 ( .A(n4758), .ZN(n4707) );
  NOR2_X4 U4560 ( .A1(n47), .A2(n5471), .ZN(n3386) );
  INV_X2 U4564 ( .A(n2384), .ZN(n1022) );
  INV_X2 U4579 ( .A(n3832), .ZN(n3031) );
  INV_X8 U4580 ( .A(a[11]), .ZN(n3793) );
  NOR2_X4 U4583 ( .A1(n4710), .A2(n2965), .ZN(n2321) );
  NAND2_X2 U4584 ( .A1(n6432), .A2(n2470), .ZN(n6619) );
  NOR2_X2 U4585 ( .A1(n4872), .A2(n1063), .ZN(n1331) );
  NAND2_X2 U4590 ( .A1(n4872), .A2(n1063), .ZN(n1330) );
  INV_X2 U4591 ( .A(n3491), .ZN(n2481) );
  NOR2_X4 U4595 ( .A1(n2536), .A2(n2535), .ZN(n1260) );
  INV_X4 U4596 ( .A(n1431), .ZN(n850) );
  NAND2_X4 U4598 ( .A1(n5887), .A2(n3476), .ZN(n5320) );
  INV_X4 U4599 ( .A(n3893), .ZN(n1486) );
  NOR2_X4 U4603 ( .A1(n6349), .A2(n3318), .ZN(n3359) );
  NAND2_X2 U4617 ( .A1(n1431), .A2(n4316), .ZN(n852) );
  NAND2_X2 U4626 ( .A1(n6628), .A2(n2696), .ZN(n6621) );
  INV_X2 U4644 ( .A(n3996), .ZN(n3997) );
  INV_X2 U4652 ( .A(n6645), .ZN(n945) );
  AOI22_X2 U4658 ( .A1(n3878), .A2(n3879), .B1(n3880), .B2(n6181), .ZN(n3881)
         );
  NAND2_X2 U4659 ( .A1(n2024), .A2(n6351), .ZN(n6622) );
  NOR2_X4 U4687 ( .A1(n1526), .A2(n1525), .ZN(n3711) );
  INV_X1 U4688 ( .A(n4637), .ZN(n2904) );
  NAND2_X2 U4689 ( .A1(n1975), .A2(n4571), .ZN(n1976) );
  NAND2_X1 U4699 ( .A1(n17), .A2(n3778), .ZN(n6625) );
  INV_X2 U4794 ( .A(n4301), .ZN(n4291) );
  INV_X1 U4796 ( .A(n3008), .ZN(n2273) );
  NAND2_X1 U4798 ( .A1(b[19]), .A2(a[1]), .ZN(n6629) );
  NAND2_X2 U4833 ( .A1(n6627), .A2(n6628), .ZN(n6630) );
  NAND2_X2 U4844 ( .A1(n6629), .A2(n6630), .ZN(n2924) );
  INV_X1 U4879 ( .A(b[19]), .ZN(n6627) );
  NAND2_X4 U4892 ( .A1(a[7]), .A2(n1287), .ZN(n4800) );
  INV_X2 U4894 ( .A(n2567), .ZN(n773) );
  NAND2_X1 U4899 ( .A1(n3616), .A2(n2567), .ZN(n774) );
  NOR3_X4 U4921 ( .A1(n3511), .A2(n4151), .A3(n5666), .ZN(n4156) );
  INV_X4 U4950 ( .A(n2349), .ZN(n1957) );
  NAND2_X1 U4976 ( .A1(n4298), .A2(n4299), .ZN(n6633) );
  NAND2_X2 U4981 ( .A1(n6633), .A2(n6634), .ZN(n2173) );
  INV_X2 U5009 ( .A(n2851), .ZN(n6058) );
  NAND2_X2 U5010 ( .A1(n4763), .A2(n3545), .ZN(n2673) );
  XNOR2_X1 U5011 ( .A(n4260), .B(n4243), .ZN(n1122) );
  INV_X1 U5015 ( .A(n4243), .ZN(n4259) );
  NOR2_X1 U5018 ( .A1(n4800), .A2(b[5]), .ZN(n6638) );
  NAND2_X1 U5020 ( .A1(n3342), .A2(n4800), .ZN(n3821) );
  OR2_X1 U5023 ( .A1(n4800), .A2(b[0]), .ZN(n986) );
  NOR3_X1 U5037 ( .A1(n5865), .A2(n5864), .A3(n5875), .ZN(n5866) );
  NAND2_X1 U5052 ( .A1(n1034), .A2(n3382), .ZN(n1814) );
  INV_X2 U5053 ( .A(n1906), .ZN(n1904) );
  INV_X2 U5066 ( .A(n4881), .ZN(n1086) );
  NAND2_X2 U5078 ( .A1(n1786), .A2(n4867), .ZN(n1563) );
  NAND2_X2 U5096 ( .A1(n669), .A2(n668), .ZN(n4867) );
  NOR2_X2 U5102 ( .A1(n6635), .A2(n6023), .ZN(\d[32] ) );
  NOR2_X4 U5131 ( .A1(n5313), .A2(n5312), .ZN(n3105) );
  NOR2_X4 U5141 ( .A1(n5851), .A2(n5854), .ZN(n5312) );
  NOR2_X2 U5157 ( .A1(n5865), .A2(n5864), .ZN(n5395) );
  NAND3_X2 U5163 ( .A1(n996), .A2(n1357), .A3(n5887), .ZN(n5865) );
  NAND2_X2 U5166 ( .A1(n1382), .A2(n6636), .ZN(n4899) );
  OAI21_X1 U5169 ( .B1(n4915), .B2(n4913), .A(n4914), .ZN(n6636) );
  AOI21_X2 U5170 ( .B1(n3491), .B2(n281), .A(n3546), .ZN(n2853) );
  NAND2_X4 U5173 ( .A1(n1849), .A2(n1009), .ZN(n3491) );
  NAND2_X2 U5191 ( .A1(n344), .A2(n6601), .ZN(n5095) );
  NAND2_X2 U5193 ( .A1(n881), .A2(n4976), .ZN(n344) );
  NAND2_X2 U5200 ( .A1(n3202), .A2(n3615), .ZN(n6257) );
  NOR3_X2 U5214 ( .A1(n1883), .A2(n6638), .A3(n6637), .ZN(n2528) );
  NAND2_X2 U5216 ( .A1(n1887), .A2(n1886), .ZN(n6637) );
  NAND3_X2 U5230 ( .A1(n1692), .A2(n2265), .A3(n1691), .ZN(n5794) );
  NOR2_X2 U5248 ( .A1(n5777), .A2(n5768), .ZN(n2265) );
  NOR2_X2 U5251 ( .A1(n3884), .A2(n3883), .ZN(n51) );
  NAND2_X2 U5253 ( .A1(n3225), .A2(n3876), .ZN(n3884) );
  NOR2_X2 U5264 ( .A1(n5020), .A2(n6462), .ZN(n4925) );
  NOR2_X2 U5271 ( .A1(n6467), .A2(n6460), .ZN(n5020) );
  NAND2_X2 U5276 ( .A1(n6639), .A2(n3707), .ZN(n2109) );
  AOI21_X2 U5284 ( .B1(n266), .B2(n3902), .A(n3746), .ZN(n3745) );
  NOR2_X2 U5287 ( .A1(n3302), .A2(n3303), .ZN(n1592) );
  NAND2_X2 U5296 ( .A1(n1156), .A2(n1157), .ZN(n3302) );
  NAND2_X2 U5298 ( .A1(n6640), .A2(n3743), .ZN(n3185) );
  NAND2_X2 U5305 ( .A1(n1246), .A2(n6641), .ZN(n2529) );
  NAND4_X1 U5306 ( .A1(n2167), .A2(n2166), .A3(n2168), .A4(n2479), .ZN(n6641)
         );
  NOR2_X4 U5309 ( .A1(n4634), .A2(n1400), .ZN(n5793) );
  NAND2_X2 U5316 ( .A1(n6062), .A2(n1902), .ZN(n496) );
  NAND3_X2 U5320 ( .A1(n6111), .A2(n2908), .A3(n6133), .ZN(n6132) );
  NAND3_X2 U5321 ( .A1(n5966), .A2(n5967), .A3(n5965), .ZN(\d[45] ) );
  NAND2_X2 U5331 ( .A1(n2879), .A2(n5604), .ZN(n2878) );
  NAND2_X2 U5332 ( .A1(n839), .A2(n838), .ZN(n1120) );
  NAND2_X2 U5340 ( .A1(n1451), .A2(n6642), .ZN(n4293) );
  NAND3_X2 U5354 ( .A1(n2436), .A2(n1454), .A3(n3987), .ZN(n6642) );
  NAND3_X1 U5359 ( .A1(n6056), .A2(n3771), .A3(n1902), .ZN(n2986) );
  NAND2_X2 U5364 ( .A1(n6643), .A2(n681), .ZN(n683) );
  INV_X2 U5372 ( .A(n1351), .ZN(n6643) );
  AOI22_X2 U5414 ( .A1(n5868), .A2(n5867), .B1(n5866), .B2(n1547), .ZN(n1351)
         );
  NAND3_X1 U5419 ( .A1(n1835), .A2(n1834), .A3(n4388), .ZN(n6644) );
  NAND3_X2 U5425 ( .A1(n4587), .A2(a[2]), .A3(b[22]), .ZN(n6645) );
  NAND2_X2 U5446 ( .A1(n6062), .A2(n1902), .ZN(n6088) );
  NAND2_X2 U5456 ( .A1(n6647), .A2(n6646), .ZN(n3545) );
  OAI21_X2 U5480 ( .B1(n1651), .B2(n2536), .A(n2535), .ZN(n6646) );
  NAND2_X2 U5485 ( .A1(n1261), .A2(n1260), .ZN(n6647) );
  OAI21_X2 U5488 ( .B1(n6056), .B2(n6055), .A(n6469), .ZN(n6057) );
  INV_X4 U5494 ( .A(n6135), .ZN(n6056) );
  NAND2_X2 U5495 ( .A1(n5604), .A2(n5863), .ZN(n6135) );
  NAND2_X2 U5502 ( .A1(n6648), .A2(n2540), .ZN(n3284) );
  NAND2_X2 U5512 ( .A1(n5473), .A2(n4598), .ZN(n6648) );
  NOR2_X2 U5530 ( .A1(n4734), .A2(n2283), .ZN(n6649) );
  NOR2_X4 U5581 ( .A1(n4547), .A2(n4546), .ZN(n6650) );
  INV_X4 U5584 ( .A(n6651), .ZN(n5919) );
  NAND2_X2 U5592 ( .A1(n5809), .A2(n3672), .ZN(n6651) );
  NAND2_X2 U5603 ( .A1(n6652), .A2(n6049), .ZN(n6061) );
  INV_X2 U5604 ( .A(n6138), .ZN(n6652) );
  NAND2_X2 U5613 ( .A1(n2452), .A2(n6275), .ZN(n2450) );
  NAND2_X2 U5629 ( .A1(n6653), .A2(n944), .ZN(n2323) );
  NAND2_X2 U5653 ( .A1(n943), .A2(n942), .ZN(n6653) );
  NAND3_X1 U5656 ( .A1(n3940), .A2(n3939), .A3(n2838), .ZN(n1414) );
  NAND2_X2 U5659 ( .A1(n4927), .A2(n4926), .ZN(n4928) );
  NAND2_X2 U5660 ( .A1(n6512), .A2(n2503), .ZN(n4927) );
  AOI22_X2 U5665 ( .A1(n216), .A2(n257), .B1(n4526), .B2(n2117), .ZN(n2166) );
  BUF_X4 U5673 ( .A(n2131), .Z(n6655) );
  NAND2_X2 U5674 ( .A1(n802), .A2(n3014), .ZN(n1070) );
  NAND3_X2 U5676 ( .A1(n1384), .A2(a[13]), .A3(a[14]), .ZN(n805) );
  INV_X8 U5678 ( .A(a[15]), .ZN(n1384) );
  INV_X2 U5681 ( .A(n6656), .ZN(n963) );
  NAND2_X2 U5685 ( .A1(n6658), .A2(n6657), .ZN(n6260) );
  INV_X2 U5686 ( .A(n3323), .ZN(n6657) );
  NAND2_X2 U5702 ( .A1(n6660), .A2(n6659), .ZN(n2301) );
  NAND2_X2 U5706 ( .A1(n5017), .A2(n5019), .ZN(n6660) );
  NOR2_X4 U5707 ( .A1(n3689), .A2(n6523), .ZN(n5928) );
  NAND2_X2 U5708 ( .A1(n2329), .A2(n6519), .ZN(n2862) );
  BUF_X4 U5714 ( .A(n5597), .Z(n6661) );
  NOR2_X2 U5727 ( .A1(n5156), .A2(n5157), .ZN(n5159) );
  NOR2_X2 U5733 ( .A1(n1379), .A2(n1378), .ZN(n5156) );
  NAND2_X2 U5734 ( .A1(n3634), .A2(n5085), .ZN(n2418) );
  NAND3_X2 U5736 ( .A1(n1830), .A2(n2050), .A3(n2051), .ZN(n6403) );
  NAND2_X2 U5755 ( .A1(n2301), .A2(n6662), .ZN(n4952) );
  NAND3_X1 U5760 ( .A1(n5017), .A2(n5019), .A3(n968), .ZN(n6662) );
  INV_X4 U5761 ( .A(n6663), .ZN(n886) );
  NOR2_X2 U5765 ( .A1(n3598), .A2(n4994), .ZN(n6664) );
  NAND2_X2 U5769 ( .A1(n6025), .A2(n2851), .ZN(n6138) );
  NAND2_X2 U5771 ( .A1(n6135), .A2(n3157), .ZN(n6025) );
  NAND2_X2 U5773 ( .A1(n2105), .A2(n2106), .ZN(n909) );
  OAI21_X2 U5775 ( .B1(n2775), .B2(n3200), .A(n4522), .ZN(n2106) );
  NAND2_X2 U5776 ( .A1(n5061), .A2(n5060), .ZN(n5130) );
  NAND2_X2 U5788 ( .A1(n273), .A2(n272), .ZN(n5061) );
  NOR2_X2 U5791 ( .A1(n6665), .A2(n1377), .ZN(n1749) );
  INV_X2 U5792 ( .A(n2756), .ZN(n6665) );
  NAND2_X2 U5796 ( .A1(n133), .A2(n3109), .ZN(n2756) );
  NAND2_X2 U5797 ( .A1(n6666), .A2(n2466), .ZN(n2464) );
  NAND2_X2 U5799 ( .A1(n4620), .A2(n2467), .ZN(n6666) );
  NAND2_X2 U5804 ( .A1(n6667), .A2(n6466), .ZN(n6675) );
  INV_X2 U5805 ( .A(n3598), .ZN(n6667) );
  OAI21_X2 U5807 ( .B1(n3199), .B2(n608), .A(n2009), .ZN(n2455) );
  AOI22_X2 U5815 ( .A1(n4495), .A2(n3187), .B1(n6212), .B2(b[20]), .ZN(n2009)
         );
  INV_X2 U5817 ( .A(n1070), .ZN(n588) );
  NAND2_X2 U5819 ( .A1(n5208), .A2(n5209), .ZN(n1506) );
  INV_X2 U5826 ( .A(n6275), .ZN(n3210) );
  OAI21_X2 U5833 ( .B1(n1651), .B2(n2536), .A(n2535), .ZN(n6275) );
  NAND2_X2 U5837 ( .A1(n2919), .A2(n4453), .ZN(n6668) );
  XNOR2_X2 U5840 ( .A(n4448), .B(n4449), .ZN(n11) );
  AOI21_X2 U5843 ( .B1(n4436), .B2(n4437), .A(n4435), .ZN(n4448) );
  NAND2_X2 U5844 ( .A1(n2296), .A2(n4382), .ZN(n3021) );
  NAND2_X2 U5851 ( .A1(n6216), .A2(n4031), .ZN(n2296) );
  AOI21_X1 U5853 ( .B1(n1013), .B2(n1902), .A(n5638), .ZN(n5640) );
  NAND2_X2 U5862 ( .A1(n4524), .A2(n4525), .ZN(n2318) );
  NAND2_X2 U5870 ( .A1(n1583), .A2(n3064), .ZN(n4525) );
  NOR2_X2 U5871 ( .A1(n6192), .A2(n639), .ZN(n6669) );
  NAND2_X2 U5872 ( .A1(n871), .A2(n872), .ZN(n6192) );
  NAND2_X4 U5879 ( .A1(n6671), .A2(n6670), .ZN(n1263) );
  NAND2_X2 U5881 ( .A1(n2511), .A2(n4497), .ZN(n6670) );
  NAND2_X2 U5884 ( .A1(n190), .A2(n189), .ZN(n6671) );
  NOR2_X2 U5885 ( .A1(n3743), .A2(n6673), .ZN(n6672) );
  INV_X2 U5886 ( .A(n3744), .ZN(n6673) );
  AOI22_X2 U5887 ( .A1(n5454), .A2(b[2]), .B1(n314), .B2(n2249), .ZN(n251) );
  NAND2_X2 U5894 ( .A1(a[15]), .A2(n2284), .ZN(n1060) );
  NOR2_X4 U5899 ( .A1(a[13]), .A2(a[14]), .ZN(n2284) );
  NAND2_X2 U5904 ( .A1(n673), .A2(n672), .ZN(n2574) );
  NAND2_X2 U5908 ( .A1(n1627), .A2(n1507), .ZN(n672) );
  INV_X4 U5910 ( .A(n6398), .ZN(n673) );
  NAND2_X2 U5918 ( .A1(n4858), .A2(n4857), .ZN(n4885) );
  NAND3_X2 U5921 ( .A1(n2640), .A2(n2639), .A3(n4856), .ZN(n4857) );
  NOR2_X2 U5924 ( .A1(n2316), .A2(n2978), .ZN(n1228) );
  NOR2_X4 U5926 ( .A1(n1989), .A2(n1987), .ZN(n2316) );
  AOI21_X2 U5928 ( .B1(n5265), .B2(n5264), .A(n5263), .ZN(n5332) );
  NAND3_X2 U5933 ( .A1(n1412), .A2(n1409), .A3(n1411), .ZN(n5265) );
  BUF_X4 U5934 ( .A(n5226), .Z(n6674) );
  NAND2_X2 U5938 ( .A1(n3299), .A2(n6675), .ZN(n5113) );
  NAND2_X2 U5941 ( .A1(n6676), .A2(n785), .ZN(n5115) );
  NAND2_X2 U5942 ( .A1(n6443), .A2(n784), .ZN(n6676) );
  OAI21_X2 U5955 ( .B1(n229), .B2(n4881), .A(n6677), .ZN(n4900) );
  NAND2_X2 U5968 ( .A1(n6214), .A2(n1041), .ZN(n6677) );
  AOI21_X2 U5977 ( .B1(n1420), .B2(n5204), .A(n6678), .ZN(n1418) );
  NOR2_X2 U5983 ( .A1(n5204), .A2(n5202), .ZN(n6678) );
  NAND3_X2 U5989 ( .A1(n6679), .A2(n1727), .A3(n6458), .ZN(n4863) );
  NOR2_X2 U5991 ( .A1(n1220), .A2(n1221), .ZN(n6679) );
  NAND2_X2 U5998 ( .A1(n6680), .A2(n6073), .ZN(n6166) );
  NAND2_X4 U6022 ( .A1(n1990), .A2(n1076), .ZN(n6092) );
  NAND2_X2 U3497 ( .A1(n1603), .A2(a[22]), .ZN(n1389) );
  INV_X4 U94 ( .A(b[0]), .ZN(n3540) );
  NOR2_X2 U1887 ( .A1(n3431), .A2(b[2]), .ZN(n3667) );
  NAND2_X2 U3604 ( .A1(n1476), .A2(n1477), .ZN(n1475) );
  NAND2_X2 U3602 ( .A1(n1475), .A2(n1473), .ZN(n4164) );
  NAND2_X2 U1230 ( .A1(n2201), .A2(n2200), .ZN(n3410) );
  INV_X2 U2906 ( .A(b[5]), .ZN(n3835) );
  INV_X2 U247 ( .A(n4802), .ZN(n6259) );
  INV_X1 U445 ( .A(n5298), .ZN(n6154) );
  INV_X2 U3358 ( .A(n3382), .ZN(n1807) );
  INV_X4 U5339 ( .A(n4305), .ZN(n3355) );
  INV_X1 U33 ( .A(n3519), .ZN(n6681) );
  NOR2_X2 U132 ( .A1(n5828), .A2(n6681), .ZN(n6189) );
  INV_X1 U179 ( .A(n3164), .ZN(n6682) );
  NOR2_X2 U264 ( .A1(n5591), .A2(n6682), .ZN(n3758) );
  INV_X1 U278 ( .A(n3164), .ZN(n6683) );
  NOR2_X2 U332 ( .A1(n5616), .A2(n6683), .ZN(n3759) );
  AND2_X2 U333 ( .A1(n5984), .A2(n5985), .ZN(n5988) );
  AOI21_X1 U335 ( .B1(n2863), .B2(n6077), .A(n6684), .ZN(n3767) );
  INV_X1 U418 ( .A(n6084), .ZN(n6684) );
  AOI21_X1 U447 ( .B1(n6077), .B2(n6078), .A(n6076), .ZN(n6084) );
  INV_X1 U473 ( .A(n6072), .ZN(n6685) );
  NOR2_X2 U517 ( .A1(n6685), .A2(n6001), .ZN(n2711) );
  INV_X1 U606 ( .A(n1615), .ZN(n6686) );
  NAND2_X2 U607 ( .A1(n6686), .A2(n1613), .ZN(n1608) );
  NAND3_X1 U608 ( .A1(n434), .A2(n3341), .A3(n432), .ZN(n995) );
  AND2_X2 U680 ( .A1(n5203), .A2(n1103), .ZN(n5205) );
  INV_X2 U697 ( .A(n5506), .ZN(n5504) );
  NAND2_X1 U819 ( .A1(n5455), .A2(n5456), .ZN(n5506) );
  OAI211_X1 U829 ( .C1(b[17]), .C2(b[16]), .A(a[23]), .B(n6687), .ZN(n5419) );
  NAND2_X1 U1024 ( .A1(b[17]), .A2(b[16]), .ZN(n6687) );
  INV_X2 U1034 ( .A(n6688), .ZN(n6634) );
  NOR2_X2 U1041 ( .A1(n4298), .A2(n4299), .ZN(n6688) );
  AND2_X2 U1077 ( .A1(n4182), .A2(n4228), .ZN(n3457) );
  OR2_X2 U1135 ( .A1(n1034), .A2(n3382), .ZN(n1806) );
  AND2_X2 U1138 ( .A1(n490), .A2(n491), .ZN(n2012) );
  NOR2_X1 U1175 ( .A1(n3575), .A2(n4919), .ZN(n951) );
  OR2_X2 U1202 ( .A1(n5303), .A2(n5298), .ZN(n4) );
  INV_X2 U1267 ( .A(n6689), .ZN(n5649) );
  NOR2_X2 U1268 ( .A1(n4135), .A2(n4136), .ZN(n6689) );
  OAI21_X1 U1281 ( .B1(n4111), .B2(n4490), .A(n4110), .ZN(n4114) );
  AND2_X2 U1395 ( .A1(n4104), .A2(n4103), .ZN(n6586) );
  INV_X2 U1599 ( .A(n1764), .ZN(n4190) );
  NAND2_X1 U1625 ( .A1(b[0]), .A2(n4933), .ZN(n1764) );
  INV_X1 U1759 ( .A(n262), .ZN(n2721) );
  NOR2_X1 U1789 ( .A1(n2748), .A2(n3888), .ZN(n262) );
  INV_X1 U1791 ( .A(n4332), .ZN(n6690) );
  OAI21_X2 U1969 ( .B1(n3730), .B2(n6690), .A(n6213), .ZN(n1004) );
  INV_X1 U1971 ( .A(n5352), .ZN(n3661) );
  AOI21_X1 U1972 ( .B1(n2570), .B2(n2568), .A(n5274), .ZN(n5352) );
  INV_X1 U2111 ( .A(n4046), .ZN(n5118) );
  NOR2_X1 U2162 ( .A1(n3639), .A2(n6188), .ZN(n4046) );
  INV_X2 U2163 ( .A(n6691), .ZN(n6626) );
  NOR2_X2 U2170 ( .A1(n17), .A2(n3778), .ZN(n6691) );
  INV_X2 U2205 ( .A(n4004), .ZN(n6692) );
  NAND2_X2 U2366 ( .A1(n6692), .A2(n4002), .ZN(n2523) );
  INV_X1 U2419 ( .A(n1171), .ZN(n2439) );
  NAND2_X1 U2455 ( .A1(n4842), .A2(n4841), .ZN(n1171) );
  INV_X1 U2467 ( .A(n940), .ZN(n2720) );
  NAND2_X1 U2481 ( .A1(n4510), .A2(n4511), .ZN(n940) );
  INV_X1 U2487 ( .A(n1189), .ZN(n5427) );
  NAND2_X1 U2517 ( .A1(b[16]), .A2(a[23]), .ZN(n1189) );
  OR2_X2 U2520 ( .A1(n401), .A2(n4802), .ZN(n599) );
  INV_X1 U2541 ( .A(n6694), .ZN(n2960) );
  NOR2_X2 U2574 ( .A1(n2965), .A2(n4710), .ZN(n6694) );
  INV_X2 U2592 ( .A(n6695), .ZN(n669) );
  NOR2_X2 U2627 ( .A1(n1785), .A2(n4865), .ZN(n6695) );
  AND2_X2 U2651 ( .A1(n4165), .A2(n4166), .ZN(n3616) );
  OR2_X2 U2659 ( .A1(n4596), .A2(n4597), .ZN(n1855) );
  INV_X1 U2660 ( .A(n6659), .ZN(n968) );
  NOR2_X1 U2664 ( .A1(n5016), .A2(n5015), .ZN(n6659) );
  INV_X2 U2725 ( .A(n6696), .ZN(n33) );
  OAI22_X1 U2766 ( .A1(n2656), .A2(b[15]), .B1(n805), .B2(n35), .ZN(n6696) );
  AOI22_X1 U2810 ( .A1(n865), .A2(n5074), .B1(b[11]), .B2(n2675), .ZN(n6446)
         );
  OR2_X2 U2812 ( .A1(n414), .A2(n4848), .ZN(n6458) );
  OR2_X2 U2835 ( .A1(n4767), .A2(b[21]), .ZN(n219) );
  AND3_X1 U2849 ( .A1(n5010), .A2(n4749), .A3(n4750), .ZN(n3281) );
  INV_X1 U2855 ( .A(n479), .ZN(n985) );
  NAND2_X1 U2868 ( .A1(a[7]), .A2(n4948), .ZN(n479) );
  INV_X1 U2877 ( .A(n5240), .ZN(n6697) );
  NAND2_X2 U2885 ( .A1(n5241), .A2(n6697), .ZN(n761) );
  OR2_X2 U2889 ( .A1(n4753), .A2(b[5]), .ZN(n4750) );
  INV_X1 U2908 ( .A(a[15]), .ZN(n2958) );
  INV_X2 U3053 ( .A(a[15]), .ZN(n2577) );
  INV_X1 U3125 ( .A(a[7]), .ZN(n6698) );
  NOR2_X2 U3322 ( .A1(n6698), .A2(b[9]), .ZN(n3880) );
  NAND2_X2 U3388 ( .A1(n4291), .A2(n3583), .ZN(n4313) );
  NAND2_X1 U3605 ( .A1(n4302), .A2(n1836), .ZN(n3583) );
  OR2_X2 U3669 ( .A1(n4543), .A2(b[4]), .ZN(n1476) );
  AND2_X2 U3872 ( .A1(b[0]), .A2(n2098), .ZN(n4514) );
  INV_X1 U3874 ( .A(a[7]), .ZN(n6699) );
  NAND2_X2 U3881 ( .A1(a[5]), .A2(n6699), .ZN(n4536) );
endmodule



    module conf_int_mul__noFF__arch_agnos__w_wrapper_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 ( 
        clk, rst, a, b, d, d__acc, acc__sel );
  input [23:0] a;
  input [23:0] b;
  output [63:0] d;
  input [63:0] d__acc;
  input clk, rst, acc__sel;
  wire   n35, n34, n37, n36, n38, n45, n30, n33, n90, n31, n42, n55, n54, n39,
         n51, n44, n43, n32, n56, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n82, n81, n80, n75, n77, n76, n85, n84, n83, n41, n40, n86, n87,
         n88, n89, n92, n91, n93, n79, n78, n1, n47, n46, n49, n48, n50, n52,
         n53, n57, n58, n59, n60, n61, n64, n94;
  wire   [47:0] d__apx;

  NAND2_X1 U96 ( .A1(n35), .A2(n34), .ZN(d[51]) );
  NAND2_X1 U141 ( .A1(n37), .A2(n36), .ZN(d[44]) );
  NAND2_X1 U142 ( .A1(n38), .A2(n45), .ZN(d[60]) );
  NAND2_X1 U143 ( .A1(n30), .A2(n33), .ZN(d[61]) );
  NAND2_X2 U144 ( .A1(d__apx[45]), .A2(n90), .ZN(n30) );
  NAND2_X1 U145 ( .A1(n31), .A2(n42), .ZN(d[47]) );
  NAND2_X1 U146 ( .A1(n55), .A2(n54), .ZN(d[48]) );
  NAND2_X1 U147 ( .A1(n39), .A2(n51), .ZN(d[50]) );
  NAND2_X1 U148 ( .A1(n44), .A2(n43), .ZN(d[56]) );
  INV_X8 U149 ( .A(acc__sel), .ZN(n90) );
  NAND2_X1 U150 ( .A1(n32), .A2(n56), .ZN(d[63]) );
  NAND2_X2 U151 ( .A1(d__apx[31]), .A2(n90), .ZN(n31) );
  NAND2_X2 U152 ( .A1(d__apx[47]), .A2(n90), .ZN(n32) );
  OAI21_X1 U154 ( .B1(d__apx[5]), .B2(acc__sel), .A(n65), .ZN(d[21]) );
  OAI21_X1 U155 ( .B1(d__apx[6]), .B2(acc__sel), .A(n66), .ZN(d[22]) );
  OAI21_X1 U156 ( .B1(d__apx[7]), .B2(acc__sel), .A(n67), .ZN(d[23]) );
  OAI21_X1 U157 ( .B1(d__apx[8]), .B2(acc__sel), .A(n68), .ZN(d[24]) );
  OAI21_X1 U158 ( .B1(d__apx[9]), .B2(acc__sel), .A(n69), .ZN(d[25]) );
  OAI21_X1 U159 ( .B1(d__apx[10]), .B2(acc__sel), .A(n70), .ZN(d[26]) );
  OAI21_X1 U160 ( .B1(d__apx[11]), .B2(acc__sel), .A(n71), .ZN(d[27]) );
  OAI21_X1 U161 ( .B1(d__apx[12]), .B2(acc__sel), .A(n72), .ZN(d[28]) );
  OAI21_X1 U162 ( .B1(d__apx[13]), .B2(acc__sel), .A(n73), .ZN(d[29]) );
  OAI21_X1 U163 ( .B1(d__apx[14]), .B2(acc__sel), .A(n74), .ZN(d[30]) );
  OAI21_X1 U164 ( .B1(d__apx[15]), .B2(acc__sel), .A(n82), .ZN(d[31]) );
  NAND2_X1 U165 ( .A1(n81), .A2(n80), .ZN(d[32]) );
  OAI21_X1 U166 ( .B1(d__apx[17]), .B2(acc__sel), .A(n75), .ZN(d[33]) );
  NAND2_X1 U167 ( .A1(n77), .A2(n76), .ZN(d[35]) );
  NAND2_X1 U168 ( .A1(n85), .A2(n84), .ZN(d[36]) );
  OAI21_X1 U169 ( .B1(d__apx[21]), .B2(acc__sel), .A(n83), .ZN(d[37]) );
  NAND2_X1 U170 ( .A1(n41), .A2(n40), .ZN(d[46]) );
  NAND2_X2 U171 ( .A1(d__apx[35]), .A2(n90), .ZN(n35) );
  NAND2_X2 U172 ( .A1(d__apx[28]), .A2(n90), .ZN(n37) );
  NAND2_X2 U173 ( .A1(d__apx[44]), .A2(n90), .ZN(n38) );
  NAND2_X2 U174 ( .A1(d__apx[34]), .A2(n90), .ZN(n39) );
  NAND2_X2 U175 ( .A1(d__apx[30]), .A2(n90), .ZN(n41) );
  OAI21_X1 U176 ( .B1(d__apx[27]), .B2(acc__sel), .A(n86), .ZN(d[43]) );
  OAI21_X1 U177 ( .B1(d__apx[23]), .B2(acc__sel), .A(n87), .ZN(d[39]) );
  OAI21_X1 U178 ( .B1(d__apx[22]), .B2(acc__sel), .A(n88), .ZN(d[38]) );
  OAI21_X1 U179 ( .B1(d__apx[24]), .B2(acc__sel), .A(n89), .ZN(d[40]) );
  NAND2_X1 U180 ( .A1(n92), .A2(n91), .ZN(d[41]) );
  OAI21_X1 U181 ( .B1(d__apx[42]), .B2(acc__sel), .A(n93), .ZN(d[58]) );
  NAND2_X1 U183 ( .A1(n79), .A2(n78), .ZN(d[34]) );
  LOGIC0_X1 U184 ( .Z(n1) );
  NAND2_X2 U185 ( .A1(d__apx[40]), .A2(n90), .ZN(n44) );
  NAND2_X2 U186 ( .A1(d__apx[43]), .A2(n90), .ZN(n47) );
  NAND2_X1 U187 ( .A1(n47), .A2(n46), .ZN(d[59]) );
  NAND2_X2 U188 ( .A1(d__apx[29]), .A2(n90), .ZN(n49) );
  NAND2_X1 U189 ( .A1(n49), .A2(n48), .ZN(d[45]) );
  OAI21_X1 U190 ( .B1(d__apx[33]), .B2(acc__sel), .A(n50), .ZN(d[49]) );
  OAI21_X1 U191 ( .B1(d__apx[46]), .B2(acc__sel), .A(n52), .ZN(d[62]) );
  OAI21_X1 U192 ( .B1(d__apx[39]), .B2(acc__sel), .A(n53), .ZN(d[55]) );
  NAND2_X2 U193 ( .A1(d__apx[32]), .A2(n90), .ZN(n55) );
  OAI21_X1 U194 ( .B1(d__apx[41]), .B2(acc__sel), .A(n57), .ZN(d[57]) );
  OAI21_X1 U195 ( .B1(d__apx[38]), .B2(acc__sel), .A(n58), .ZN(d[54]) );
  OAI21_X1 U196 ( .B1(d__apx[37]), .B2(acc__sel), .A(n59), .ZN(d[53]) );
  OAI21_X1 U197 ( .B1(d__apx[26]), .B2(acc__sel), .A(n60), .ZN(d[42]) );
  OAI21_X1 U198 ( .B1(d__apx[36]), .B2(acc__sel), .A(n61), .ZN(d[52]) );
  OAI21_X1 U199 ( .B1(d__apx[4]), .B2(acc__sel), .A(n64), .ZN(d[20]) );
  NAND2_X2 U200 ( .A1(d__apx[19]), .A2(n90), .ZN(n77) );
  NAND2_X2 U201 ( .A1(d__apx[18]), .A2(n90), .ZN(n79) );
  NAND2_X2 U202 ( .A1(d__apx[16]), .A2(n90), .ZN(n81) );
  NAND2_X2 U203 ( .A1(d__apx[25]), .A2(n90), .ZN(n92) );
  AND2_X1 U204 ( .A1(acc__sel), .A2(d__acc[0]), .ZN(d[0]) );
  AND2_X1 U205 ( .A1(acc__sel), .A2(d__acc[1]), .ZN(d[1]) );
  AND2_X1 U206 ( .A1(acc__sel), .A2(d__acc[2]), .ZN(d[2]) );
  AND2_X1 U207 ( .A1(acc__sel), .A2(d__acc[3]), .ZN(d[3]) );
  AND2_X1 U208 ( .A1(acc__sel), .A2(d__acc[4]), .ZN(d[4]) );
  AND2_X1 U209 ( .A1(acc__sel), .A2(d__acc[5]), .ZN(d[5]) );
  AND2_X1 U210 ( .A1(acc__sel), .A2(d__acc[6]), .ZN(d[6]) );
  AND2_X1 U211 ( .A1(acc__sel), .A2(d__acc[7]), .ZN(d[7]) );
  AND2_X1 U212 ( .A1(acc__sel), .A2(d__acc[8]), .ZN(d[8]) );
  AND2_X1 U213 ( .A1(acc__sel), .A2(d__acc[9]), .ZN(d[9]) );
  AND2_X1 U214 ( .A1(acc__sel), .A2(d__acc[10]), .ZN(d[10]) );
  AND2_X1 U215 ( .A1(acc__sel), .A2(d__acc[11]), .ZN(d[11]) );
  AND2_X1 U216 ( .A1(acc__sel), .A2(d__acc[12]), .ZN(d[12]) );
  AND2_X1 U217 ( .A1(acc__sel), .A2(d__acc[13]), .ZN(d[13]) );
  AND2_X1 U218 ( .A1(acc__sel), .A2(d__acc[14]), .ZN(d[14]) );
  AND2_X1 U219 ( .A1(acc__sel), .A2(d__acc[15]), .ZN(d[15]) );
  MUX2_X1 U220 ( .A(d__apx[0]), .B(d__acc[16]), .S(acc__sel), .Z(d[16]) );
  NAND2_X2 U118 ( .A1(acc__sel), .A2(d__acc[49]), .ZN(n50) );
  NAND2_X2 U99 ( .A1(acc__sel), .A2(d__acc[40]), .ZN(n89) );
  NAND2_X2 U106 ( .A1(acc__sel), .A2(d__acc[54]), .ZN(n58) );
  NAND2_X2 U104 ( .A1(acc__sel), .A2(d__acc[38]), .ZN(n88) );
  NAND2_X2 U101 ( .A1(acc__sel), .A2(d__acc[39]), .ZN(n87) );
  NAND2_X2 U110 ( .A1(acc__sel), .A2(d__acc[52]), .ZN(n61) );
  NAND2_X2 U114 ( .A1(acc__sel), .A2(d__acc[58]), .ZN(n93) );
  NAND2_X2 U107 ( .A1(acc__sel), .A2(d__acc[55]), .ZN(n53) );
  NAND2_X2 U121 ( .A1(acc__sel), .A2(d__acc[62]), .ZN(n52) );
  NAND2_X2 U126 ( .A1(acc__sel), .A2(d__acc[43]), .ZN(n86) );
  NAND2_X2 U109 ( .A1(acc__sel), .A2(d__acc[53]), .ZN(n59) );
  NAND2_X2 U139 ( .A1(acc__sel), .A2(d__acc[33]), .ZN(n75) );
  NAND2_X2 U136 ( .A1(acc__sel), .A2(d__acc[31]), .ZN(n82) );
  NAND2_X2 U133 ( .A1(acc__sel), .A2(d__acc[30]), .ZN(n74) );
  NAND2_X2 U135 ( .A1(acc__sel), .A2(d__acc[29]), .ZN(n73) );
  NAND2_X2 U100 ( .A1(acc__sel), .A2(d__acc[28]), .ZN(n72) );
  NAND2_X2 U138 ( .A1(acc__sel), .A2(d__acc[37]), .ZN(n83) );
  conf_int_mul__noFF__arch_agnos_OP_BITWIDTH22_DATA_PATH_BITWIDTH24 mul__inst ( 
        .clk(clk), .rst(n1), .a(a), .b(b), .\d[47] (d__apx[47]), .\d[44] (
        d__apx[44]), .\d[43] (d__apx[43]), .\d[40] (d__apx[40]), .\d[37]_BAR (
        d__apx[37]), .\d[34] (d__apx[34]), .\d[31] (d__apx[31]), .\d[28] (
        d__apx[28]), .\d[16] (d__apx[16]), .\d[1] (d__apx[1]), .\d[0] (
        d__apx[0]), .\d[33]_BAR (d__apx[33]), .\d[27]_BAR (d__apx[27]), 
        .\d[26]_BAR (d__apx[26]), .\d[24]_BAR (d__apx[24]), .\d[23]_BAR (
        d__apx[23]), .\d[21]_BAR (d__apx[21]), .\d[15]_BAR (d__apx[15]), 
        .\d[14]_BAR (d__apx[14]), .\d[11]_BAR (d__apx[11]), .\d[9]_BAR (
        d__apx[9]), .\d[6]_BAR (d__apx[6]), .\d[4]_BAR (d__apx[4]), 
        .\d[42]_BAR (d__apx[42]), .\d[41]_BAR (d__apx[41]), .\d[30] (
        d__apx[30]), .\d[22]_BAR (d__apx[22]), .\d[46]_BAR (d__apx[46]), 
        .\d[35] (d__apx[35]), .\d[19] (d__apx[19]), .\d[10]_BAR (d__apx[10]), 
        .\d[8]_BAR (d__apx[8]), .\d[5]_BAR (d__apx[5]), .\d[3] (d__apx[3]), 
        .\d[29] (d__apx[29]), .\d[7]_BAR (d__apx[7]), .\d[32] (d__apx[32]), 
        .\d[39]_BAR (d__apx[39]), .\d[12]_BAR (d__apx[12]), .\d[2] (d__apx[2]), 
        .\d[36]_BAR (d__apx[36]), .\d[25] (d__apx[25]), .\d[13]_BAR (
        d__apx[13]), .\d[38]_BAR (d__apx[38]), .\d[20] (d__apx[20]), .\d[18] (
        d__apx[18]), .\d[45] (d__apx[45]), .\d[17]_BAR (d__apx[17]) );
  NAND2_X2 U108 ( .A1(acc__sel), .A2(d__acc[63]), .ZN(n56) );
  NAND2_X2 U95 ( .A1(acc__sel), .A2(d__acc[20]), .ZN(n64) );
  NAND2_X2 U122 ( .A1(acc__sel), .A2(d__acc[21]), .ZN(n65) );
  NAND2_X2 U102 ( .A1(acc__sel), .A2(d__acc[22]), .ZN(n66) );
  NAND2_X2 U105 ( .A1(acc__sel), .A2(d__acc[23]), .ZN(n67) );
  NAND2_X2 U137 ( .A1(acc__sel), .A2(d__acc[24]), .ZN(n68) );
  NAND2_X2 U129 ( .A1(acc__sel), .A2(d__acc[25]), .ZN(n69) );
  NAND2_X2 U113 ( .A1(acc__sel), .A2(d__acc[51]), .ZN(n34) );
  NAND2_X2 U97 ( .A1(acc__sel), .A2(d__acc[41]), .ZN(n91) );
  NAND2_X2 U128 ( .A1(acc__sel), .A2(d__acc[35]), .ZN(n76) );
  NAND2_X2 U111 ( .A1(acc__sel), .A2(d__acc[56]), .ZN(n43) );
  NAND2_X2 U130 ( .A1(acc__sel), .A2(d__acc[32]), .ZN(n80) );
  NAND2_X2 U116 ( .A1(acc__sel), .A2(d__acc[59]), .ZN(n46) );
  NAND2_X2 U140 ( .A1(acc__sel), .A2(d__acc[36]), .ZN(n84) );
  NAND2_X2 U117 ( .A1(acc__sel), .A2(d__acc[60]), .ZN(n45) );
  NAND2_X2 U119 ( .A1(acc__sel), .A2(d__acc[61]), .ZN(n33) );
  NAND2_X2 U134 ( .A1(acc__sel), .A2(d__acc[34]), .ZN(n78) );
  NAND2_X2 U124 ( .A1(acc__sel), .A2(d__acc[45]), .ZN(n48) );
  NAND2_X2 U115 ( .A1(acc__sel), .A2(d__acc[50]), .ZN(n51) );
  NAND2_X2 U125 ( .A1(acc__sel), .A2(d__acc[44]), .ZN(n36) );
  NAND2_X2 U120 ( .A1(acc__sel), .A2(d__acc[48]), .ZN(n54) );
  NAND2_X2 U127 ( .A1(acc__sel), .A2(d__acc[46]), .ZN(n40) );
  NAND2_X2 U123 ( .A1(acc__sel), .A2(d__acc[47]), .ZN(n42) );
  MUX2_X2 U221 ( .A(d__apx[1]), .B(d__acc[17]), .S(acc__sel), .Z(d[17]) );
  MUX2_X2 U94 ( .A(d__apx[2]), .B(d__acc[18]), .S(acc__sel), .Z(d[18]) );
  NAND2_X2 U93 ( .A1(d__apx[20]), .A2(n90), .ZN(n85) );
  NAND2_X2 U98 ( .A1(acc__sel), .A2(d__acc[42]), .ZN(n60) );
  NAND2_X2 U112 ( .A1(acc__sel), .A2(d__acc[57]), .ZN(n57) );
  NAND2_X2 U131 ( .A1(acc__sel), .A2(d__acc[27]), .ZN(n71) );
  NAND2_X2 U132 ( .A1(acc__sel), .A2(d__acc[26]), .ZN(n70) );
  INV_X1 U103 ( .A(n94), .ZN(d[19]) );
  AOI22_X1 U153 ( .A1(d__acc[19]), .A2(acc__sel), .B1(n90), .B2(d__apx[3]), 
        .ZN(n94) );
endmodule

