library verilog;
use verilog.vl_types.all;
entity AOI21_X2_func is
    port(
        A               : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        ZN              : out    vl_logic
    );
end AOI21_X2_func;
