module conf_int_mul__noFF__arch_agnos_OP_BITWIDTH18_DATA_PATH_BITWIDTH26 ( clk, 
        racc, rapx, a, b, \d[24] , \d[23] , \d[22] , \d[20] , \d[19] , \d[17] , 
        \d[9] , \d[1] , \d[0] , \d[16]_BAR , \d[4]_BAR , \d[2]_BAR , 
        \d[15]_BAR , \d[14] , \d[18] , \d[21] , \d[10] , \d[6] , \d[5] , 
        \d[13] , \d[12] , \d[3] , \d[11]_BAR , \d[8] , \d[7]  );
  input [25:0] a;
  input [14:0] b;
  input clk, racc, rapx;
  output \d[24] , \d[23] , \d[22] , \d[20] , \d[19] , \d[17] , \d[9] , \d[1] ,
         \d[0] , \d[16]_BAR , \d[4]_BAR , \d[2]_BAR , \d[15]_BAR , \d[14] ,
         \d[18] , \d[21] , \d[10] , \d[6] , \d[5] , \d[13] , \d[12] , \d[3] ,
         \d[11]_BAR , \d[8] , \d[7] ;
  wire   \intadd_0/SUM[2] , n1, n2, n3, n6, n8, n9, n10, n11, n13, n14, n16,
         n17, n18, n19, n20, n22, n23, n25, n27, n29, n30, n31, n32, n35, n36,
         n37, n38, n40, n41, n42, n44, n45, n46, n47, n50, n51, n52, n53, n55,
         n56, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97, n98, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n126, n127, n128, n129, n130, n131, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n155, n156, n157, n158, n159,
         n160, n161, n163, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n200, n201, n202, n203, n204, n205, n206, n207, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n224, n225, n226, n227, n228, n229, n230, n231, n233, n234,
         n235, n236, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n250, n253, n254, n255, n256, n257, n259, n260, n261,
         n262, n263, n264, n265, n268, n269, n270, n271, n272, n273, n274,
         n277, n278, n281, n282, n283, n285, n286, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n321, n322, n325, n326, n327, n328, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n342, n343,
         n344, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n361, n362, n363, n364, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n382, n383, n384, n385,
         n387, n388, n389, n390, n391, n392, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n404, n405, n406, n407, n411, n412, n416,
         n417, n418, n420, n422, n427, n428, n429, n431, n432, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n452, n453, n454, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n511, n512, n513, n514, n515, n516, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n571, n572, n573, n574, n575, n576, n578, n579, n580, n583, n584,
         n587, n589, n590, n591, n592, n593, n596, n597, n598, n599, n600,
         n601, n602, n603, n605, n606, n608, n610, n612, n613, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n652, n653, n654, n655, n656, n657, n658, n659, n661, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n682, n683, n684, n685, n686, n687,
         n689, n691, n692, n693, n694, n695, n696, n697, n698, n700, n701,
         n703, n704, n705, n706, n707, n708, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n737, n738,
         n741, n742, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n775, n776, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n826, n827, n828, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n923, n924, n925,
         n926, n927, n928, n929, n930, n932, n933, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n954, n955, n956, n957, n959, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n973, n974, n975,
         n976, n977, n978, n979, n982, n983, n984, n986, n987, n988, n989,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1036, n1038, n1039, n1040, n1042, n1043, n1045, n1046, n1047,
         n1048, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1104, n1105, n1107, n1108, n1109, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1172, n1173, n1174,
         n1175, n1176, n1177, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1202, n1203, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1225, n1226, n1227, n1228,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1239, n1241,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1291, n1292, n1293, n1294, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1314, n1315, n1316, n1317,
         n1318, n1319, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1339,
         n1340, n1342, n1343, n1344, n1345, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1359, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1452, n1453, n1454, n1455, n1456, n1457, n1459, n1461, n1463,
         n1464, n1465, n1466, n1467, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1484, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1502, n1503, n1504, n1505, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1515, n1517, n1518, n1519, n1520, n1521, n1522,
         n1525, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1536,
         n1537, n1538, n1539, n1540, n1545, n1547, n1550, n1551, n1552, n1553,
         n1554, n1555, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1577, n1578, n1579, n1580, n1585, n1586, n1587, n1588, n1589, n1591,
         n1593, n1594, n1595, n1596, n1597, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1643, n1644, n1645, n1646, n1647,
         n1649, n1650, n1651, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765;
  assign \d[7]  = \intadd_0/SUM[2] ;

  BUF_X4 U3 ( .A(n1390), .Z(n27) );
  NOR2_X2 U6 ( .A1(n600), .A2(n1395), .ZN(n133) );
  NAND2_X2 U7 ( .A1(n391), .A2(n390), .ZN(n838) );
  INV_X1 U8 ( .A(n1114), .ZN(n30) );
  INV_X2 U9 ( .A(n1505), .ZN(n794) );
  NOR2_X2 U11 ( .A1(n802), .A2(a[8]), .ZN(n1221) );
  NOR2_X2 U12 ( .A1(n845), .A2(n40), .ZN(n856) );
  INV_X4 U15 ( .A(n1410), .ZN(n38) );
  INV_X1 U19 ( .A(n606), .ZN(n50) );
  INV_X1 U20 ( .A(n1364), .ZN(n319) );
  NAND2_X2 U33 ( .A1(n127), .A2(n1), .ZN(n186) );
  INV_X2 U34 ( .A(n2), .ZN(n1) );
  NOR2_X2 U36 ( .A1(n3), .A2(n116), .ZN(n933) );
  NAND2_X2 U37 ( .A1(n932), .A2(n1663), .ZN(n3) );
  NAND2_X2 U43 ( .A1(n484), .A2(n1427), .ZN(n483) );
  NAND3_X2 U44 ( .A1(n1278), .A2(n1277), .A3(n1424), .ZN(n1427) );
  INV_X4 U45 ( .A(n444), .ZN(n178) );
  INV_X4 U48 ( .A(n109), .ZN(n108) );
  INV_X4 U50 ( .A(n1328), .ZN(n885) );
  NAND2_X2 U54 ( .A1(n6), .A2(n1272), .ZN(n1423) );
  INV_X2 U55 ( .A(n272), .ZN(n6) );
  NAND2_X2 U56 ( .A1(n1268), .A2(n1267), .ZN(n272) );
  NAND2_X2 U57 ( .A1(n84), .A2(n179), .ZN(n1128) );
  NOR2_X2 U62 ( .A1(n1423), .A2(n486), .ZN(n485) );
  NAND2_X2 U63 ( .A1(n715), .A2(n714), .ZN(n73) );
  NAND2_X2 U64 ( .A1(n1521), .A2(n513), .ZN(n714) );
  INV_X4 U65 ( .A(n1683), .ZN(n805) );
  INV_X4 U66 ( .A(n881), .ZN(n737) );
  XNOR2_X2 U70 ( .A(n1235), .B(n1234), .ZN(n446) );
  NAND2_X2 U71 ( .A1(n670), .A2(n669), .ZN(n1234) );
  NAND2_X2 U72 ( .A1(n84), .A2(n1750), .ZN(n1255) );
  NAND2_X2 U74 ( .A1(n11), .A2(n10), .ZN(n9) );
  BUF_X2 U90 ( .A(n307), .Z(n13) );
  NOR2_X2 U91 ( .A1(n1646), .A2(n14), .ZN(n913) );
  NAND2_X2 U92 ( .A1(n411), .A2(n597), .ZN(n14) );
  NAND2_X2 U97 ( .A1(n771), .A2(n213), .ZN(n212) );
  NAND2_X2 U106 ( .A1(b[14]), .A2(n1683), .ZN(n18) );
  NAND3_X2 U108 ( .A1(n1608), .A2(n1188), .A3(n90), .ZN(n85) );
  NAND2_X2 U109 ( .A1(n146), .A2(n1197), .ZN(n327) );
  NAND2_X2 U110 ( .A1(n19), .A2(n319), .ZN(n314) );
  NOR3_X2 U111 ( .A1(n359), .A2(n1363), .A3(n600), .ZN(n19) );
  NAND2_X2 U115 ( .A1(n623), .A2(n685), .ZN(n110) );
  NAND2_X4 U116 ( .A1(n745), .A2(n547), .ZN(n685) );
  AOI21_X2 U119 ( .B1(n1046), .B2(b[8]), .A(n1045), .ZN(n1050) );
  NAND2_X2 U122 ( .A1(n36), .A2(n204), .ZN(n197) );
  XNOR2_X1 U125 ( .A(n808), .B(n1125), .ZN(n1122) );
  XNOR2_X1 U126 ( .A(n805), .B(n1512), .ZN(n1028) );
  NAND2_X1 U128 ( .A1(n179), .A2(a[20]), .ZN(n1067) );
  NAND2_X1 U132 ( .A1(n273), .A2(n1596), .ZN(n761) );
  NAND3_X1 U138 ( .A1(n1315), .A2(n1314), .A3(n376), .ZN(\d[8] ) );
  BUF_X4 U141 ( .A(n1496), .Z(n25) );
  INV_X4 U142 ( .A(n1221), .ZN(n29) );
  INV_X4 U146 ( .A(n1164), .ZN(n55) );
  OR2_X2 U151 ( .A1(n1235), .A2(n29), .ZN(n1217) );
  INV_X4 U154 ( .A(n257), .ZN(n160) );
  AND2_X4 U155 ( .A1(n1188), .A2(n951), .ZN(n31) );
  NOR2_X4 U162 ( .A1(n300), .A2(n306), .ZN(n1086) );
  NAND2_X2 U164 ( .A1(n734), .A2(n1645), .ZN(n331) );
  AND2_X4 U165 ( .A1(n1333), .A2(n1400), .ZN(n36) );
  NAND3_X1 U168 ( .A1(n1167), .A2(n1083), .A3(n1709), .ZN(n373) );
  NAND2_X1 U169 ( .A1(n41), .A2(n159), .ZN(n1391) );
  OR2_X1 U170 ( .A1(n1453), .A2(n1452), .ZN(n957) );
  INV_X1 U172 ( .A(n661), .ZN(n627) );
  INV_X2 U173 ( .A(n1400), .ZN(n37) );
  INV_X2 U174 ( .A(n352), .ZN(n1189) );
  INV_X2 U176 ( .A(n1306), .ZN(n51) );
  NAND2_X1 U177 ( .A1(n575), .A2(n574), .ZN(n573) );
  INV_X4 U178 ( .A(n1160), .ZN(n40) );
  INV_X4 U179 ( .A(a[12]), .ZN(n991) );
  INV_X2 U181 ( .A(a[14]), .ZN(n1001) );
  OR2_X2 U184 ( .A1(n1325), .A2(n1328), .ZN(n549) );
  NAND2_X1 U185 ( .A1(n377), .A2(n957), .ZN(n1315) );
  XNOR2_X1 U188 ( .A(n1422), .B(n1421), .ZN(\intadd_0/SUM[2] ) );
  XOR2_X1 U190 ( .A(n627), .B(n705), .Z(n959) );
  NOR2_X2 U191 ( .A1(n1399), .A2(n1086), .ZN(n1316) );
  INV_X4 U192 ( .A(n1616), .ZN(n41) );
  INV_X4 U193 ( .A(n719), .ZN(n42) );
  INV_X1 U194 ( .A(n1459), .ZN(n898) );
  NAND2_X2 U198 ( .A1(n480), .A2(n481), .ZN(n1192) );
  INV_X2 U200 ( .A(n1149), .ZN(n644) );
  INV_X1 U201 ( .A(n1384), .ZN(n45) );
  XNOR2_X1 U202 ( .A(n1378), .B(n1377), .ZN(n1380) );
  BUF_X4 U205 ( .A(n1291), .Z(n561) );
  INV_X2 U207 ( .A(n1291), .ZN(n1200) );
  OR2_X2 U208 ( .A1(n1112), .A2(n1113), .ZN(n599) );
  INV_X4 U210 ( .A(n1177), .ZN(n46) );
  INV_X1 U216 ( .A(n1249), .ZN(n1244) );
  NAND2_X2 U218 ( .A1(n402), .A2(n1658), .ZN(n849) );
  INV_X2 U221 ( .A(n1136), .ZN(n52) );
  NAND2_X2 U222 ( .A1(n810), .A2(n811), .ZN(n525) );
  NAND2_X2 U224 ( .A1(n1027), .A2(n1026), .ZN(n779) );
  INV_X2 U230 ( .A(a[9]), .ZN(n994) );
  INV_X2 U231 ( .A(a[13]), .ZN(n695) );
  INV_X4 U232 ( .A(n991), .ZN(n53) );
  INV_X1 U235 ( .A(a[23]), .ZN(n946) );
  INV_X1 U236 ( .A(a[22]), .ZN(n840) );
  NAND2_X1 U238 ( .A1(n57), .A2(n769), .ZN(n56) );
  BUF_X4 U239 ( .A(n1074), .Z(n57) );
  INV_X4 U242 ( .A(n235), .ZN(n233) );
  INV_X4 U244 ( .A(n394), .ZN(n1270) );
  NOR2_X2 U248 ( .A1(n845), .A2(n1140), .ZN(n894) );
  NAND3_X2 U249 ( .A1(n1444), .A2(n1441), .A3(n1424), .ZN(n1279) );
  NAND2_X2 U251 ( .A1(n71), .A2(n69), .ZN(n400) );
  NAND2_X2 U252 ( .A1(n59), .A2(n1316), .ZN(n1317) );
  NAND3_X1 U256 ( .A1(n870), .A2(n1108), .A3(n871), .ZN(n61) );
  NAND2_X2 U257 ( .A1(n60), .A2(n61), .ZN(n441) );
  NAND2_X2 U258 ( .A1(n264), .A2(n692), .ZN(n60) );
  INV_X2 U259 ( .A(n1098), .ZN(n230) );
  INV_X2 U261 ( .A(n64), .ZN(n63) );
  NOR2_X2 U262 ( .A1(n1043), .A2(n1065), .ZN(n64) );
  INV_X4 U263 ( .A(n769), .ZN(n1153) );
  NAND2_X1 U267 ( .A1(n1160), .A2(n65), .ZN(n527) );
  INV_X4 U277 ( .A(n72), .ZN(n715) );
  NAND2_X2 U279 ( .A1(n73), .A2(n1220), .ZN(n554) );
  AOI21_X2 U280 ( .B1(n1722), .B2(n242), .A(n1292), .ZN(n1220) );
  NAND3_X2 U284 ( .A1(n1528), .A2(n95), .A3(n96), .ZN(n243) );
  NAND2_X2 U285 ( .A1(n94), .A2(n1289), .ZN(n244) );
  NAND2_X2 U287 ( .A1(n552), .A2(n832), .ZN(n74) );
  NAND2_X2 U289 ( .A1(n809), .A2(n941), .ZN(n917) );
  NOR2_X4 U291 ( .A1(n318), .A2(n1366), .ZN(n809) );
  NAND2_X4 U293 ( .A1(n584), .A2(n583), .ZN(n626) );
  NOR2_X2 U294 ( .A1(n798), .A2(a[24]), .ZN(n1137) );
  NOR2_X2 U296 ( .A1(n813), .A2(n814), .ZN(n1194) );
  NOR2_X2 U297 ( .A1(n1064), .A2(n1063), .ZN(n813) );
  INV_X4 U298 ( .A(n753), .ZN(n399) );
  NOR2_X4 U299 ( .A1(n798), .A2(n1164), .ZN(n1071) );
  AND2_X4 U302 ( .A1(n618), .A2(b[8]), .ZN(n948) );
  NOR2_X4 U305 ( .A1(n1607), .A2(n752), .ZN(n621) );
  NAND2_X2 U306 ( .A1(n1058), .A2(n757), .ZN(n1059) );
  NAND2_X2 U308 ( .A1(n812), .A2(n1091), .ZN(n1092) );
  BUF_X4 U312 ( .A(n1033), .Z(n77) );
  OAI21_X2 U313 ( .B1(n993), .B2(n1410), .A(n1508), .ZN(n225) );
  NAND2_X2 U317 ( .A1(n770), .A2(n1098), .ZN(n871) );
  NAND2_X2 U319 ( .A1(n79), .A2(n78), .ZN(n896) );
  NAND2_X2 U323 ( .A1(n80), .A2(n612), .ZN(n790) );
  NAND2_X4 U327 ( .A1(n1257), .A2(n1510), .ZN(n143) );
  NAND2_X2 U329 ( .A1(n845), .A2(n53), .ZN(n893) );
  NAND2_X4 U332 ( .A1(n81), .A2(n1059), .ZN(n1188) );
  NAND2_X2 U333 ( .A1(n145), .A2(n1057), .ZN(n81) );
  NAND2_X2 U336 ( .A1(n311), .A2(n1247), .ZN(n308) );
  NAND2_X2 U338 ( .A1(n282), .A2(n283), .ZN(n82) );
  INV_X4 U340 ( .A(n1509), .ZN(n496) );
  BUF_X4 U341 ( .A(n84), .Z(n83) );
  INV_X8 U344 ( .A(n995), .ZN(n84) );
  INV_X4 U345 ( .A(n1197), .ZN(n654) );
  NOR2_X1 U349 ( .A1(n394), .A2(a[24]), .ZN(n217) );
  NAND2_X1 U350 ( .A1(n40), .A2(n394), .ZN(n857) );
  NAND2_X2 U352 ( .A1(n91), .A2(n253), .ZN(n1243) );
  NAND3_X2 U356 ( .A1(n93), .A2(n472), .A3(n901), .ZN(n1136) );
  NAND2_X2 U359 ( .A1(n95), .A2(n96), .ZN(n94) );
  INV_X4 U363 ( .A(n747), .ZN(n97) );
  NAND2_X2 U367 ( .A1(n101), .A2(n100), .ZN(n907) );
  NAND2_X2 U368 ( .A1(n877), .A2(n639), .ZN(n100) );
  NAND2_X2 U370 ( .A1(n707), .A2(n858), .ZN(n102) );
  NAND2_X2 U371 ( .A1(n757), .A2(n967), .ZN(n858) );
  NAND2_X2 U372 ( .A1(n966), .A2(n841), .ZN(n954) );
  NOR2_X2 U375 ( .A1(n103), .A2(n314), .ZN(n318) );
  INV_X8 U376 ( .A(n104), .ZN(n257) );
  NAND3_X2 U379 ( .A1(n106), .A2(n1232), .A3(n105), .ZN(n242) );
  NAND2_X2 U380 ( .A1(n1216), .A2(n29), .ZN(n105) );
  NOR2_X2 U381 ( .A1(n545), .A2(n555), .ZN(n1232) );
  NAND2_X2 U382 ( .A1(n1211), .A2(n1235), .ZN(n106) );
  NAND2_X4 U383 ( .A1(n107), .A2(n108), .ZN(n1065) );
  NAND2_X2 U387 ( .A1(n111), .A2(n725), .ZN(n623) );
  NAND2_X2 U388 ( .A1(n149), .A2(n150), .ZN(n111) );
  NAND2_X4 U389 ( .A1(n114), .A2(n112), .ZN(n330) );
  INV_X4 U390 ( .A(n113), .ZN(n112) );
  NAND2_X2 U391 ( .A1(n726), .A2(n725), .ZN(n113) );
  INV_X4 U392 ( .A(n685), .ZN(n114) );
  NOR2_X2 U394 ( .A1(n622), .A2(n621), .ZN(n766) );
  NAND2_X2 U395 ( .A1(n116), .A2(n44), .ZN(n292) );
  INV_X4 U396 ( .A(n1630), .ZN(n116) );
  NAND2_X1 U402 ( .A1(n1001), .A2(n120), .ZN(n119) );
  BUF_X4 U403 ( .A(n468), .Z(n121) );
  NAND2_X4 U405 ( .A1(n468), .A2(n808), .ZN(n412) );
  AOI21_X1 U407 ( .B1(n928), .B2(n468), .A(n689), .ZN(n1063) );
  NAND2_X2 U412 ( .A1(n1021), .A2(n263), .ZN(n724) );
  NAND2_X2 U413 ( .A1(n123), .A2(n1029), .ZN(n1111) );
  NAND2_X2 U414 ( .A1(n282), .A2(n57), .ZN(n123) );
  NAND2_X2 U415 ( .A1(n257), .A2(a[19]), .ZN(n1077) );
  INV_X4 U417 ( .A(n1021), .ZN(n723) );
  NAND2_X2 U418 ( .A1(n781), .A2(n552), .ZN(n1484) );
  NAND2_X4 U428 ( .A1(n126), .A2(n218), .ZN(n1176) );
  NAND2_X2 U429 ( .A1(n220), .A2(n221), .ZN(n126) );
  NOR2_X2 U431 ( .A1(n188), .A2(n187), .ZN(n127) );
  AOI21_X2 U433 ( .B1(n1130), .B2(n1239), .A(n805), .ZN(n1003) );
  NAND2_X2 U436 ( .A1(n1520), .A2(n1200), .ZN(n128) );
  NAND2_X2 U437 ( .A1(n793), .A2(n986), .ZN(n713) );
  XNOR2_X2 U443 ( .A(n808), .B(n928), .ZN(n1075) );
  NOR2_X2 U445 ( .A1(n293), .A2(n129), .ZN(\d[23] ) );
  NAND2_X2 U447 ( .A1(n131), .A2(n130), .ZN(n784) );
  INV_X2 U449 ( .A(n477), .ZN(n131) );
  NAND2_X2 U451 ( .A1(n247), .A2(a[19]), .ZN(n1057) );
  NOR2_X2 U456 ( .A1(n1188), .A2(n951), .ZN(n363) );
  NAND2_X2 U457 ( .A1(n1647), .A2(n727), .ZN(n729) );
  NAND2_X2 U462 ( .A1(n628), .A2(n1356), .ZN(n910) );
  NAND2_X2 U470 ( .A1(n1222), .A2(n1221), .ZN(n1211) );
  INV_X8 U473 ( .A(n1053), .ZN(n489) );
  NAND2_X4 U474 ( .A1(n489), .A2(n682), .ZN(n684) );
  BUF_X4 U475 ( .A(n888), .Z(n138) );
  NAND3_X2 U476 ( .A1(n139), .A2(n152), .A3(n1350), .ZN(\d[21] ) );
  NAND2_X2 U479 ( .A1(n141), .A2(n140), .ZN(n516) );
  INV_X2 U480 ( .A(n1643), .ZN(n140) );
  INV_X2 U481 ( .A(n1018), .ZN(n141) );
  INV_X4 U488 ( .A(n1379), .ZN(n1332) );
  NAND2_X2 U490 ( .A1(n304), .A2(n854), .ZN(n303) );
  INV_X4 U499 ( .A(n1538), .ZN(n150) );
  INV_X8 U500 ( .A(n143), .ZN(n845) );
  NAND2_X2 U501 ( .A1(n144), .A2(n666), .ZN(\d[11]_BAR ) );
  NAND2_X2 U502 ( .A1(n664), .A2(n665), .ZN(n144) );
  NAND2_X2 U504 ( .A1(n336), .A2(a[15]), .ZN(n1027) );
  NAND2_X2 U511 ( .A1(n979), .A2(n1410), .ZN(n982) );
  NAND2_X2 U513 ( .A1(n1249), .A2(n1756), .ZN(n710) );
  NAND2_X2 U523 ( .A1(n917), .A2(n1369), .ZN(n148) );
  INV_X2 U524 ( .A(n1487), .ZN(n1469) );
  NAND2_X1 U525 ( .A1(n1621), .A2(n512), .ZN(n613) );
  AOI21_X2 U526 ( .B1(n176), .B2(n1020), .A(n442), .ZN(n512) );
  NAND2_X2 U528 ( .A1(n1270), .A2(n57), .ZN(n1007) );
  NOR2_X4 U531 ( .A1(n203), .A2(n1072), .ZN(n1179) );
  NAND3_X2 U536 ( .A1(n418), .A2(n153), .A3(n330), .ZN(n417) );
  NAND2_X2 U539 ( .A1(n1336), .A2(n1337), .ZN(n1348) );
  NAND3_X2 U540 ( .A1(n654), .A2(n1619), .A3(n678), .ZN(n155) );
  NAND2_X2 U543 ( .A1(n1518), .A2(n156), .ZN(n444) );
  XNOR2_X2 U546 ( .A(n1174), .B(n1173), .ZN(n867) );
  NAND2_X2 U548 ( .A1(n160), .A2(a[11]), .ZN(n906) );
  NAND2_X2 U551 ( .A1(n1743), .A2(n1528), .ZN(n161) );
  NAND2_X2 U553 ( .A1(n1034), .A2(n1538), .ZN(n725) );
  NAND2_X2 U559 ( .A1(n166), .A2(n461), .ZN(n169) );
  NAND2_X2 U562 ( .A1(n172), .A2(n170), .ZN(n930) );
  INV_X2 U564 ( .A(n246), .ZN(n171) );
  OAI21_X2 U565 ( .B1(n173), .B2(n246), .A(n1115), .ZN(n172) );
  NAND2_X2 U568 ( .A1(n1332), .A2(n175), .ZN(n712) );
  NOR2_X2 U571 ( .A1(n1352), .A2(n1627), .ZN(n844) );
  NAND2_X2 U572 ( .A1(n1555), .A2(n443), .ZN(n656) );
  NAND2_X2 U573 ( .A1(n179), .A2(a[15]), .ZN(n963) );
  NAND2_X1 U574 ( .A1(n179), .A2(a[10]), .ZN(n1256) );
  NOR2_X1 U576 ( .A1(n179), .A2(n55), .ZN(n216) );
  NAND2_X2 U580 ( .A1(n1157), .A2(n1156), .ZN(n181) );
  NAND2_X2 U583 ( .A1(n186), .A2(n184), .ZN(n183) );
  NAND2_X2 U586 ( .A1(n1540), .A2(n1336), .ZN(n185) );
  NOR2_X2 U587 ( .A1(n631), .A2(n1496), .ZN(n187) );
  NAND2_X4 U588 ( .A1(n661), .A2(n1294), .ZN(n1496) );
  NAND3_X2 U591 ( .A1(n193), .A2(n190), .A3(n1319), .ZN(n189) );
  NOR2_X2 U592 ( .A1(n191), .A2(n1385), .ZN(n190) );
  NAND2_X2 U593 ( .A1(n1219), .A2(n192), .ZN(n191) );
  NOR2_X2 U594 ( .A1(n631), .A2(n1616), .ZN(n192) );
  NAND3_X2 U595 ( .A1(n316), .A2(n315), .A3(n1311), .ZN(n628) );
  AOI21_X2 U597 ( .B1(n195), .B2(n427), .A(n431), .ZN(n194) );
  NOR2_X2 U598 ( .A1(n197), .A2(n196), .ZN(n195) );
  INV_X2 U600 ( .A(n432), .ZN(n198) );
  INV_X2 U604 ( .A(n1367), .ZN(n1294) );
  NAND2_X2 U605 ( .A1(n201), .A2(n200), .ZN(n1367) );
  AOI22_X1 U608 ( .A1(n1188), .A2(n1168), .B1(n1189), .B2(n951), .ZN(n202) );
  NOR2_X4 U609 ( .A1(n1070), .A2(n1071), .ZN(n203) );
  OR2_X2 U610 ( .A1(n783), .A2(n205), .ZN(n390) );
  NAND2_X2 U611 ( .A1(n783), .A2(n205), .ZN(n392) );
  INV_X2 U612 ( .A(n77), .ZN(n205) );
  NAND2_X2 U613 ( .A1(n207), .A2(n206), .ZN(n783) );
  NAND2_X1 U614 ( .A1(n1623), .A2(n877), .ZN(n206) );
  INV_X4 U618 ( .A(n210), .ZN(n986) );
  NAND2_X2 U622 ( .A1(a[17]), .A2(n948), .ZN(n976) );
  NAND2_X2 U623 ( .A1(n22), .A2(n460), .ZN(n977) );
  NAND2_X2 U624 ( .A1(n792), .A2(n791), .ZN(n210) );
  AOI22_X2 U625 ( .A1(n559), .A2(n1678), .B1(n212), .B2(n157), .ZN(n1368) );
  NOR2_X4 U626 ( .A1(n1176), .A2(n676), .ZN(n1177) );
  NAND3_X2 U627 ( .A1(n180), .A2(n215), .A3(n214), .ZN(n676) );
  NOR2_X2 U629 ( .A1(n217), .A2(n216), .ZN(n215) );
  NAND2_X1 U631 ( .A1(n412), .A2(n40), .ZN(n219) );
  NAND2_X2 U632 ( .A1(n467), .A2(n1054), .ZN(n220) );
  NAND2_X2 U638 ( .A1(n556), .A2(n387), .ZN(n888) );
  NAND2_X2 U639 ( .A1(n225), .A2(n1227), .ZN(n1202) );
  NAND2_X2 U642 ( .A1(n1412), .A2(n1022), .ZN(n224) );
  NAND2_X2 U643 ( .A1(n901), .A2(n988), .ZN(n226) );
  NAND2_X2 U645 ( .A1(n987), .A2(n848), .ZN(n235) );
  NAND3_X2 U650 ( .A1(n240), .A2(n238), .A3(n244), .ZN(n787) );
  NOR2_X2 U651 ( .A1(n239), .A2(n1233), .ZN(n238) );
  NAND2_X2 U653 ( .A1(n242), .A2(n241), .ZN(n240) );
  AOI21_X2 U657 ( .B1(n1052), .B2(n1114), .A(n1113), .ZN(n1115) );
  NOR2_X2 U658 ( .A1(n914), .A2(n1051), .ZN(n1113) );
  NOR2_X2 U660 ( .A1(n264), .A2(n265), .ZN(n246) );
  NAND2_X2 U661 ( .A1(n871), .A2(n870), .ZN(n264) );
  NAND2_X2 U663 ( .A1(n247), .A2(a[8]), .ZN(n1253) );
  INV_X4 U664 ( .A(n1131), .ZN(n247) );
  NAND2_X2 U667 ( .A1(n915), .A2(n271), .ZN(n1261) );
  NAND2_X2 U668 ( .A1(n313), .A2(n916), .ZN(n902) );
  NOR2_X2 U670 ( .A1(n1439), .A2(n1438), .ZN(n487) );
  NAND2_X2 U671 ( .A1(n1439), .A2(n1438), .ZN(n488) );
  BUF_X4 U673 ( .A(n989), .Z(n253) );
  NOR2_X2 U677 ( .A1(n388), .A2(n746), .ZN(n254) );
  NOR2_X2 U680 ( .A1(n1287), .A2(n1291), .ZN(n388) );
  NAND2_X2 U681 ( .A1(n561), .A2(n1521), .ZN(n389) );
  NAND2_X2 U682 ( .A1(n819), .A2(n818), .ZN(n256) );
  NOR2_X2 U683 ( .A1(n261), .A2(n259), .ZN(n803) );
  NAND2_X2 U684 ( .A1(n260), .A2(n1457), .ZN(n259) );
  NAND2_X2 U686 ( .A1(n1030), .A2(n838), .ZN(n260) );
  NAND2_X4 U690 ( .A1(n1504), .A2(n945), .ZN(n262) );
  OAI22_X2 U692 ( .A1(n1004), .A2(n1065), .B1(n1003), .B2(n1002), .ZN(n263) );
  XNOR2_X1 U696 ( .A(n1575), .B(n1440), .ZN(\d[5] ) );
  NOR3_X2 U697 ( .A1(n485), .A2(n482), .A3(n483), .ZN(n269) );
  NOR2_X1 U698 ( .A1(n1722), .A2(n242), .ZN(n1392) );
  NAND3_X2 U700 ( .A1(n270), .A2(n1230), .A3(n242), .ZN(n786) );
  NAND2_X2 U701 ( .A1(n1258), .A2(n841), .ZN(n271) );
  NAND2_X2 U702 ( .A1(n272), .A2(n1269), .ZN(n366) );
  NAND2_X2 U703 ( .A1(n1125), .A2(n273), .ZN(n1069) );
  NAND2_X2 U704 ( .A1(n952), .A2(n273), .ZN(n886) );
  NAND2_X1 U706 ( .A1(n928), .A2(n273), .ZN(n574) );
  INV_X8 U708 ( .A(n776), .ZN(n273) );
  NAND2_X1 U709 ( .A1(n274), .A2(n1416), .ZN(n1417) );
  NOR2_X4 U710 ( .A1(n1416), .A2(n274), .ZN(n566) );
  NAND2_X2 U711 ( .A1(n565), .A2(n1414), .ZN(n274) );
  NAND3_X2 U714 ( .A1(n742), .A2(n569), .A3(n567), .ZN(n277) );
  NAND2_X2 U719 ( .A1(n729), .A2(n728), .ZN(n437) );
  NAND2_X2 U720 ( .A1(n1631), .A2(n1105), .ZN(n728) );
  BUF_X4 U722 ( .A(n995), .Z(n282) );
  INV_X2 U729 ( .A(n1399), .ZN(n286) );
  NOR2_X4 U730 ( .A1(n288), .A2(n1606), .ZN(n1399) );
  NAND2_X2 U732 ( .A1(n289), .A2(n1680), .ZN(n1291) );
  NAND2_X2 U733 ( .A1(n290), .A2(n578), .ZN(n289) );
  INV_X2 U734 ( .A(n793), .ZN(n290) );
  NAND2_X1 U735 ( .A1(n299), .A2(n1630), .ZN(n291) );
  NAND2_X2 U738 ( .A1(n297), .A2(n344), .ZN(n295) );
  NOR2_X2 U740 ( .A1(n1389), .A2(n1660), .ZN(n297) );
  AOI22_X2 U744 ( .A1(n680), .A2(n857), .B1(n855), .B2(n1067), .ZN(n854) );
  NAND2_X2 U746 ( .A1(n606), .A2(n473), .ZN(n305) );
  NAND2_X2 U747 ( .A1(n1090), .A2(n1089), .ZN(n473) );
  AOI22_X2 U748 ( .A1(n326), .A2(n325), .B1(n1084), .B2(n1085), .ZN(n306) );
  NAND2_X2 U749 ( .A1(n1669), .A2(n698), .ZN(n344) );
  NAND2_X2 U757 ( .A1(n1252), .A2(n1253), .ZN(n313) );
  NAND2_X2 U759 ( .A1(n1394), .A2(n1392), .ZN(n315) );
  NOR2_X2 U761 ( .A1(n1119), .A2(n748), .ZN(n1285) );
  NOR2_X2 U765 ( .A1(n638), .A2(n2), .ZN(n321) );
  NAND2_X2 U768 ( .A1(n328), .A2(n590), .ZN(n325) );
  NAND2_X2 U769 ( .A1(n1709), .A2(n520), .ZN(n328) );
  NAND3_X2 U771 ( .A1(n331), .A2(n333), .A3(n332), .ZN(n1389) );
  NOR2_X2 U773 ( .A1(n334), .A2(n719), .ZN(n333) );
  INV_X1 U774 ( .A(n1333), .ZN(n334) );
  NAND2_X1 U776 ( .A1(n1164), .A2(n336), .ZN(n1120) );
  NAND2_X2 U778 ( .A1(n694), .A2(n693), .ZN(n497) );
  NAND2_X2 U779 ( .A1(n337), .A2(n343), .ZN(n693) );
  NAND2_X2 U781 ( .A1(n342), .A2(n671), .ZN(n694) );
  NOR2_X2 U782 ( .A1(n338), .A2(n1682), .ZN(n671) );
  INV_X2 U783 ( .A(n864), .ZN(n338) );
  NAND2_X2 U784 ( .A1(n339), .A2(n906), .ZN(n864) );
  AOI21_X2 U787 ( .B1(n1342), .B2(n344), .A(n1339), .ZN(n1340) );
  NAND2_X2 U797 ( .A1(n257), .A2(n1160), .ZN(n354) );
  NOR2_X4 U799 ( .A1(n1082), .A2(n1056), .ZN(n951) );
  AOI22_X2 U800 ( .A1(n382), .A2(n350), .B1(n1074), .B2(n732), .ZN(n1056) );
  AOI22_X2 U801 ( .A1(n355), .A2(n38), .B1(n1055), .B2(n1054), .ZN(n1082) );
  XNOR2_X2 U803 ( .A(n1511), .B(n946), .ZN(n355) );
  INV_X2 U805 ( .A(n1196), .ZN(n357) );
  AOI21_X2 U806 ( .B1(n1195), .B2(n473), .A(n358), .ZN(n1196) );
  NOR2_X2 U807 ( .A1(n50), .A2(n1193), .ZN(n358) );
  INV_X2 U808 ( .A(n1709), .ZN(n1193) );
  NAND2_X2 U811 ( .A1(n368), .A2(n364), .ZN(n367) );
  INV_X2 U816 ( .A(n364), .ZN(n361) );
  NAND2_X2 U817 ( .A1(n363), .A2(n364), .ZN(n362) );
  NAND2_X2 U819 ( .A1(n1279), .A2(n366), .ZN(n482) );
  NAND2_X1 U820 ( .A1(n366), .A2(n1423), .ZN(n1426) );
  INV_X2 U823 ( .A(n369), .ZN(n716) );
  NAND2_X2 U824 ( .A1(n369), .A2(n518), .ZN(n1157) );
  AOI21_X2 U825 ( .B1(n370), .B2(n42), .A(n1322), .ZN(n1323) );
  NAND2_X2 U826 ( .A1(n1496), .A2(n1365), .ZN(n370) );
  NAND2_X2 U827 ( .A1(n626), .A2(n1390), .ZN(n1365) );
  INV_X2 U828 ( .A(n1368), .ZN(n661) );
  NAND2_X2 U831 ( .A1(n646), .A2(n645), .ZN(n371) );
  NAND2_X2 U832 ( .A1(n643), .A2(n644), .ZN(n646) );
  INV_X2 U833 ( .A(n1301), .ZN(n372) );
  OAI21_X2 U834 ( .B1(n476), .B2(n475), .A(n474), .ZN(n1301) );
  INV_X2 U837 ( .A(n375), .ZN(n374) );
  NAND2_X1 U838 ( .A1(n1312), .A2(n23), .ZN(n376) );
  INV_X1 U839 ( .A(n1312), .ZN(n377) );
  NOR2_X2 U840 ( .A1(n378), .A2(n1453), .ZN(n1456) );
  NOR2_X2 U841 ( .A1(n1312), .A2(n1452), .ZN(n378) );
  NOR2_X4 U842 ( .A1(n379), .A2(n1611), .ZN(n1312) );
  INV_X2 U847 ( .A(n57), .ZN(n382) );
  NAND3_X2 U849 ( .A1(n29), .A2(n1207), .A3(n1208), .ZN(n383) );
  NAND2_X2 U850 ( .A1(n385), .A2(n1221), .ZN(n384) );
  NAND2_X2 U851 ( .A1(n1207), .A2(n1208), .ZN(n385) );
  NAND2_X2 U852 ( .A1(n1203), .A2(n757), .ZN(n1208) );
  AOI22_X2 U854 ( .A1(n975), .A2(n757), .B1(n974), .B2(n973), .ZN(n848) );
  NAND2_X2 U855 ( .A1(n689), .A2(a[13]), .ZN(n970) );
  NAND2_X4 U856 ( .A1(n42), .A2(n41), .ZN(n663) );
  NAND2_X2 U859 ( .A1(n1032), .A2(n392), .ZN(n391) );
  NAND2_X2 U861 ( .A1(n397), .A2(n395), .ZN(n481) );
  NOR2_X2 U863 ( .A1(n896), .A2(n396), .ZN(n795) );
  NAND2_X2 U865 ( .A1(n399), .A2(n398), .ZN(n397) );
  OAI21_X2 U869 ( .B1(n850), .B2(n849), .A(n401), .ZN(n1018) );
  NAND2_X2 U874 ( .A1(n650), .A2(n649), .ZN(n404) );
  NAND2_X2 U876 ( .A1(n593), .A2(n592), .ZN(n405) );
  BUF_X4 U877 ( .A(n1184), .Z(n406) );
  NAND2_X2 U879 ( .A1(n8), .A2(n1296), .ZN(n407) );
  NAND2_X2 U887 ( .A1(n412), .A2(n1047), .ZN(n1026) );
  NAND2_X1 U888 ( .A1(n412), .A2(n1140), .ZN(n673) );
  NAND2_X1 U889 ( .A1(n412), .A2(n55), .ZN(n1121) );
  NOR2_X2 U893 ( .A1(n417), .A2(n416), .ZN(n897) );
  NOR2_X2 U894 ( .A1(n1031), .A2(n783), .ZN(n416) );
  INV_X2 U898 ( .A(n708), .ZN(n1249) );
  OAI211_X1 U899 ( .C1(a[13]), .C2(n798), .A(n420), .B(n761), .ZN(n708) );
  NOR2_X2 U903 ( .A1(n1685), .A2(n428), .ZN(n422) );
  NAND2_X2 U907 ( .A1(n42), .A2(n1664), .ZN(n428) );
  INV_X2 U910 ( .A(n1308), .ZN(n431) );
  NOR2_X4 U911 ( .A1(n731), .A2(n750), .ZN(n1403) );
  NAND2_X2 U913 ( .A1(n439), .A2(n438), .ZN(n748) );
  NAND3_X2 U918 ( .A1(n436), .A2(n598), .A3(n599), .ZN(n440) );
  NAND2_X2 U919 ( .A1(n1119), .A2(n748), .ZN(n747) );
  NAND2_X2 U921 ( .A1(n441), .A2(n440), .ZN(n439) );
  XNOR2_X2 U922 ( .A(n1033), .B(n675), .ZN(n443) );
  NOR2_X1 U923 ( .A1(n1016), .A2(n1018), .ZN(n442) );
  NAND2_X2 U925 ( .A1(n448), .A2(n446), .ZN(n616) );
  NAND2_X2 U927 ( .A1(n659), .A2(n658), .ZN(n448) );
  INV_X4 U928 ( .A(n1241), .ZN(n1055) );
  NAND2_X2 U929 ( .A1(n452), .A2(n449), .ZN(n1213) );
  NAND2_X2 U930 ( .A1(n450), .A2(n1022), .ZN(n449) );
  NAND2_X2 U932 ( .A1(n453), .A2(n1569), .ZN(n452) );
  NOR2_X2 U933 ( .A1(a[10]), .A2(n808), .ZN(n453) );
  NOR2_X4 U940 ( .A1(n460), .A2(n459), .ZN(n591) );
  NAND2_X2 U942 ( .A1(n462), .A2(n32), .ZN(n1149) );
  NAND2_X2 U943 ( .A1(n463), .A2(n1183), .ZN(n462) );
  NAND2_X2 U944 ( .A1(n466), .A2(n737), .ZN(n463) );
  NAND2_X2 U946 ( .A1(n717), .A2(n716), .ZN(n465) );
  INV_X2 U947 ( .A(n826), .ZN(n466) );
  XNOR2_X2 U948 ( .A(n1148), .B(n519), .ZN(n1151) );
  INV_X1 U949 ( .A(n471), .ZN(n1303) );
  NAND2_X2 U950 ( .A1(n470), .A2(n469), .ZN(n1133) );
  NAND2_X2 U951 ( .A1(n52), .A2(n1164), .ZN(n469) );
  NAND2_X2 U952 ( .A1(n1152), .A2(n55), .ZN(n470) );
  NAND2_X2 U955 ( .A1(n1092), .A2(n473), .ZN(n1105) );
  NAND2_X2 U957 ( .A1(n1146), .A2(n46), .ZN(n474) );
  NOR2_X2 U958 ( .A1(n46), .A2(n1146), .ZN(n475) );
  NOR2_X2 U961 ( .A1(n785), .A2(n1148), .ZN(n477) );
  NAND2_X2 U962 ( .A1(n479), .A2(n478), .ZN(n785) );
  NAND2_X2 U963 ( .A1(n1150), .A2(n519), .ZN(n478) );
  NAND2_X2 U964 ( .A1(n608), .A2(n518), .ZN(n479) );
  AOI21_X2 U967 ( .B1(n1267), .B2(n1272), .A(n1266), .ZN(n1438) );
  NAND2_X2 U968 ( .A1(n603), .A2(n489), .ZN(n672) );
  NAND2_X2 U970 ( .A1(n936), .A2(n935), .ZN(n1072) );
  NAND2_X2 U971 ( .A1(n490), .A2(n492), .ZN(n1268) );
  NOR3_X2 U972 ( .A1(n1265), .A2(n283), .A3(n121), .ZN(n492) );
  NAND2_X2 U973 ( .A1(n1264), .A2(n846), .ZN(n490) );
  NAND3_X2 U974 ( .A1(n491), .A2(n846), .A3(n1264), .ZN(n1267) );
  INV_X2 U975 ( .A(n492), .ZN(n491) );
  AOI22_X2 U977 ( .A1(n1012), .A2(b[8]), .B1(n928), .B2(n1055), .ZN(n944) );
  NOR2_X4 U979 ( .A1(n496), .A2(n53), .ZN(n815) );
  NAND2_X2 U981 ( .A1(n497), .A2(n501), .ZN(n500) );
  NAND3_X2 U983 ( .A1(n499), .A2(n694), .A3(n693), .ZN(n498) );
  INV_X4 U984 ( .A(n502), .ZN(n1420) );
  NAND2_X2 U985 ( .A1(n502), .A2(n1436), .ZN(n1281) );
  INV_X1 U987 ( .A(n625), .ZN(n505) );
  INV_X2 U988 ( .A(n1594), .ZN(n506) );
  NAND2_X2 U989 ( .A1(n506), .A2(n697), .ZN(n507) );
  NOR2_X2 U992 ( .A1(n1681), .A2(n1008), .ZN(n675) );
  NAND2_X2 U993 ( .A1(n827), .A2(n828), .ZN(n1008) );
  BUF_X4 U999 ( .A(n1627), .Z(n511) );
  XNOR2_X1 U1000 ( .A(n1353), .B(n511), .ZN(n1354) );
  XNOR2_X2 U1001 ( .A(n1019), .B(n1623), .ZN(n818) );
  AOI21_X2 U1002 ( .B1(n572), .B2(n571), .A(n1021), .ZN(n1019) );
  NAND2_X2 U1003 ( .A1(n516), .A2(n515), .ZN(n819) );
  INV_X2 U1007 ( .A(n518), .ZN(n519) );
  INV_X4 U1009 ( .A(n1088), .ZN(n520) );
  NAND2_X2 U1012 ( .A1(n522), .A2(n755), .ZN(n521) );
  NAND3_X2 U1015 ( .A1(n460), .A2(a[18]), .A3(b[10]), .ZN(n524) );
  NAND2_X4 U1016 ( .A1(n525), .A2(n1073), .ZN(n1089) );
  NAND2_X2 U1018 ( .A1(n526), .A2(n1227), .ZN(n601) );
  OAI21_X2 U1019 ( .B1(n993), .B2(n1410), .A(n1508), .ZN(n526) );
  NAND2_X2 U1023 ( .A1(n532), .A2(n1182), .ZN(n593) );
  NOR2_X2 U1030 ( .A1(n637), .A2(n1228), .ZN(n536) );
  NAND2_X2 U1032 ( .A1(n637), .A2(n1228), .ZN(n538) );
  INV_X1 U1036 ( .A(n541), .ZN(n542) );
  NOR2_X2 U1037 ( .A1(n820), .A2(a[15]), .ZN(n1048) );
  NOR2_X4 U1040 ( .A1(n1668), .A2(n1048), .ZN(n752) );
  NAND2_X2 U1042 ( .A1(n822), .A2(n807), .ZN(n691) );
  NAND2_X2 U1044 ( .A1(n648), .A2(n46), .ZN(n650) );
  INV_X4 U1046 ( .A(a[18]), .ZN(n928) );
  XNOR2_X1 U1047 ( .A(n1370), .B(n1371), .ZN(n1304) );
  NAND3_X1 U1049 ( .A1(n283), .A2(n1412), .A3(b[8]), .ZN(n1414) );
  NAND2_X1 U1051 ( .A1(n732), .A2(n991), .ZN(n575) );
  NOR2_X1 U1052 ( .A1(n1376), .A2(n991), .ZN(n926) );
  NAND2_X1 U1054 ( .A1(n1510), .A2(n682), .ZN(n642) );
  INV_X1 U1056 ( .A(n1248), .ZN(n1245) );
  NAND2_X1 U1057 ( .A1(n1249), .A2(n1248), .ZN(n1246) );
  NOR2_X1 U1059 ( .A1(n283), .A2(n1410), .ZN(\d[0] ) );
  NOR2_X1 U1061 ( .A1(n1362), .A2(n1646), .ZN(n1359) );
  XNOR2_X1 U1062 ( .A(n250), .B(n1438), .ZN(n1440) );
  XNOR2_X1 U1063 ( .A(n1432), .B(n1431), .ZN(\d[4]_BAR ) );
  XNOR2_X1 U1064 ( .A(n1426), .B(n1428), .ZN(n1432) );
  INV_X1 U1065 ( .A(n597), .ZN(n1454) );
  NAND3_X1 U1066 ( .A1(n1312), .A2(n1311), .A3(n610), .ZN(n1314) );
  NAND2_X1 U1067 ( .A1(n1444), .A2(n1417), .ZN(\d[2]_BAR ) );
  NAND2_X2 U1068 ( .A1(n1139), .A2(n672), .ZN(n1173) );
  INV_X1 U1069 ( .A(a[20]), .ZN(n801) );
  INV_X1 U1070 ( .A(n1111), .ZN(n1112) );
  NOR2_X1 U1072 ( .A1(n1263), .A2(n928), .ZN(n927) );
  INV_X1 U1074 ( .A(n587), .ZN(n1084) );
  NAND2_X1 U1075 ( .A1(n1022), .A2(n1239), .ZN(n1023) );
  INV_X1 U1077 ( .A(n1370), .ZN(n1372) );
  INV_X1 U1078 ( .A(n1404), .ZN(n925) );
  NAND2_X2 U1080 ( .A1(n978), .A2(n1055), .ZN(n1264) );
  OAI21_X1 U1081 ( .B1(n1382), .B2(n45), .A(n1380), .ZN(n1386) );
  INV_X2 U1086 ( .A(n411), .ZN(n1453) );
  INV_X1 U1089 ( .A(n1427), .ZN(n1429) );
  XNOR2_X1 U1091 ( .A(n1443), .B(n1449), .ZN(n1445) );
  NAND2_X1 U1096 ( .A1(n1442), .A2(n1441), .ZN(n1446) );
  INV_X1 U1098 ( .A(n1433), .ZN(n1435) );
  NAND3_X1 U1099 ( .A1(n1415), .A2(n1414), .A3(n1413), .ZN(\d[1] ) );
  NOR2_X1 U1100 ( .A1(n1412), .A2(n701), .ZN(n1411) );
  XOR2_X1 U1104 ( .A(n626), .B(n27), .Z(n548) );
  INV_X4 U1106 ( .A(n1090), .ZN(n812) );
  INV_X1 U1107 ( .A(n1235), .ZN(n1223) );
  INV_X4 U1108 ( .A(n1182), .ZN(n1146) );
  AOI21_X2 U1109 ( .B1(n552), .B2(n1401), .A(n1492), .ZN(n1493) );
  NAND2_X2 U1110 ( .A1(n787), .A2(n786), .ZN(n553) );
  NOR2_X1 U1111 ( .A1(n1212), .A2(n1213), .ZN(n555) );
  BUF_X4 U1114 ( .A(n765), .Z(n558) );
  NAND2_X2 U1116 ( .A1(n771), .A2(n1186), .ZN(n560) );
  NAND2_X2 U1117 ( .A1(n564), .A2(n563), .ZN(n562) );
  NAND2_X2 U1118 ( .A1(n947), .A2(a[10]), .ZN(n564) );
  NAND2_X2 U1119 ( .A1(n568), .A2(n115), .ZN(n567) );
  NOR2_X2 U1121 ( .A1(n926), .A2(n927), .ZN(n571) );
  NAND2_X4 U1123 ( .A1(n760), .A2(n779), .ZN(n914) );
  INV_X4 U1124 ( .A(b[9]), .ZN(n618) );
  NOR2_X2 U1125 ( .A1(a[20]), .A2(n1609), .ZN(n1045) );
  AOI22_X2 U1126 ( .A1(n824), .A2(b[8]), .B1(n822), .B2(n1055), .ZN(n576) );
  NAND2_X2 U1132 ( .A1(n579), .A2(n580), .ZN(n1215) );
  NOR2_X1 U1136 ( .A1(n1425), .A2(n1424), .ZN(n1428) );
  INV_X1 U1142 ( .A(n1447), .ZN(n1448) );
  NAND2_X1 U1144 ( .A1(n823), .A2(n821), .ZN(n589) );
  NAND2_X1 U1146 ( .A1(n1088), .A2(n1193), .ZN(n590) );
  NAND2_X1 U1147 ( .A1(n368), .A2(n1167), .ZN(n1168) );
  INV_X4 U1148 ( .A(n1263), .ZN(n947) );
  NAND2_X2 U1152 ( .A1(n1254), .A2(n757), .ZN(n916) );
  NAND2_X2 U1159 ( .A1(n886), .A2(n672), .ZN(n1138) );
  NAND2_X2 U1162 ( .A1(n622), .A2(n621), .ZN(n874) );
  NOR2_X2 U1163 ( .A1(n814), .A2(n813), .ZN(n606) );
  INV_X2 U1164 ( .A(n1150), .ZN(n608) );
  NAND2_X1 U1166 ( .A1(n786), .A2(n787), .ZN(n610) );
  NAND2_X2 U1167 ( .A1(n1649), .A2(n1196), .ZN(n1198) );
  INV_X1 U1168 ( .A(n1174), .ZN(n1144) );
  NOR2_X4 U1170 ( .A1(n897), .A2(n869), .ZN(n1117) );
  NAND2_X1 U1175 ( .A1(n965), .A2(b[9]), .ZN(n619) );
  NAND2_X2 U1176 ( .A1(n605), .A2(n1283), .ZN(n1418) );
  NAND2_X1 U1180 ( .A1(n1404), .A2(n1730), .ZN(n1405) );
  NAND2_X2 U1182 ( .A1(n657), .A2(n47), .ZN(n659) );
  NAND2_X1 U1184 ( .A1(n1014), .A2(n545), .ZN(n1015) );
  INV_X4 U1186 ( .A(n951), .ZN(n1167) );
  NAND2_X1 U1189 ( .A1(n978), .A2(n820), .ZN(n791) );
  NAND2_X1 U1190 ( .A1(n867), .A2(n1175), .ZN(n633) );
  NAND2_X2 U1191 ( .A1(n632), .A2(n1172), .ZN(n634) );
  INV_X2 U1192 ( .A(n867), .ZN(n632) );
  NAND2_X1 U1195 ( .A1(n257), .A2(n1060), .ZN(n827) );
  AND2_X4 U1198 ( .A1(n1055), .A2(n994), .ZN(n1271) );
  NAND2_X1 U1199 ( .A1(n672), .A2(n1139), .ZN(n635) );
  INV_X1 U1200 ( .A(n1464), .ZN(n1465) );
  NOR2_X2 U1201 ( .A1(n1496), .A2(n631), .ZN(n638) );
  NAND2_X1 U1202 ( .A1(n955), .A2(n954), .ZN(n640) );
  NAND2_X2 U1204 ( .A1(n641), .A2(n642), .ZN(n966) );
  NAND2_X2 U1206 ( .A1(n645), .A2(n646), .ZN(n1147) );
  INV_X2 U1207 ( .A(n784), .ZN(n643) );
  NAND2_X2 U1208 ( .A1(n1166), .A2(n1165), .ZN(n647) );
  NAND2_X1 U1209 ( .A1(n1219), .A2(n25), .ZN(n1369) );
  NOR2_X2 U1210 ( .A1(n865), .A2(n1177), .ZN(n1185) );
  NAND2_X1 U1211 ( .A1(n1183), .A2(n1177), .ZN(n649) );
  INV_X1 U1212 ( .A(n1227), .ZN(n668) );
  NAND2_X2 U1214 ( .A1(n701), .A2(n1047), .ZN(n653) );
  NOR2_X4 U1216 ( .A1(n944), .A2(n943), .ZN(n1051) );
  INV_X4 U1218 ( .A(n1236), .ZN(n657) );
  INV_X2 U1221 ( .A(n896), .ZN(n1166) );
  NAND2_X1 U1222 ( .A1(n908), .A2(n1354), .ZN(n666) );
  INV_X2 U1223 ( .A(n908), .ZN(n664) );
  NAND2_X2 U1225 ( .A1(n667), .A2(n668), .ZN(n670) );
  NAND2_X1 U1227 ( .A1(n1251), .A2(n816), .ZN(n1248) );
  NAND2_X1 U1230 ( .A1(n1373), .A2(n1372), .ZN(n1374) );
  OAI21_X1 U1231 ( .B1(n1373), .B2(n1372), .A(n1371), .ZN(n1375) );
  NAND2_X1 U1232 ( .A1(n472), .A2(n901), .ZN(n1302) );
  NAND2_X1 U1234 ( .A1(n1074), .A2(n1511), .ZN(n979) );
  INV_X2 U1242 ( .A(n751), .ZN(n682) );
  INV_X1 U1243 ( .A(a[16]), .ZN(n751) );
  NOR2_X1 U1246 ( .A1(n1502), .A2(n1611), .ZN(n1422) );
  NOR2_X2 U1248 ( .A1(n605), .A2(n1283), .ZN(n1309) );
  INV_X4 U1250 ( .A(n887), .ZN(n841) );
  NOR2_X2 U1251 ( .A1(n1134), .A2(n887), .ZN(n1135) );
  NAND2_X4 U1253 ( .A1(n1181), .A2(n1180), .ZN(n1186) );
  INV_X1 U1255 ( .A(n804), .ZN(n698) );
  NAND2_X2 U1257 ( .A1(n47), .A2(n1235), .ZN(n700) );
  NAND2_X2 U1259 ( .A1(n701), .A2(n1160), .ZN(n703) );
  NAND2_X4 U1261 ( .A1(n1053), .A2(n38), .ZN(n776) );
  INV_X4 U1262 ( .A(n989), .ZN(n807) );
  NAND2_X2 U1263 ( .A1(n1491), .A2(n767), .ZN(n1492) );
  NOR2_X1 U1264 ( .A1(n1323), .A2(n1328), .ZN(n1326) );
  INV_X1 U1265 ( .A(n635), .ZN(n1143) );
  NAND2_X1 U1266 ( .A1(n635), .A2(n1174), .ZN(n1145) );
  NAND2_X2 U1268 ( .A1(n1185), .A2(n1184), .ZN(n771) );
  NAND2_X1 U1271 ( .A1(n708), .A2(n1522), .ZN(n711) );
  BUF_X4 U1273 ( .A(n968), .Z(n756) );
  NAND2_X1 U1275 ( .A1(a[18]), .A2(n845), .ZN(n778) );
  NAND2_X1 U1276 ( .A1(a[18]), .A2(n937), .ZN(n936) );
  NAND3_X2 U1277 ( .A1(n1487), .A2(n1488), .A3(n733), .ZN(n1489) );
  INV_X1 U1278 ( .A(n1185), .ZN(n1187) );
  OAI22_X1 U1280 ( .A1(n1307), .A2(n542), .B1(n1306), .B2(n1373), .ZN(n1384)
         );
  NAND2_X1 U1281 ( .A1(a[19]), .A2(n937), .ZN(n823) );
  NAND2_X2 U1282 ( .A1(n1218), .A2(n775), .ZN(n1324) );
  NAND2_X2 U1284 ( .A1(n150), .A2(n149), .ZN(n726) );
  INV_X1 U1285 ( .A(n767), .ZN(n730) );
  NAND2_X1 U1286 ( .A1(n1151), .A2(n1150), .ZN(n919) );
  NAND2_X2 U1291 ( .A1(n1504), .A2(n945), .ZN(n734) );
  INV_X1 U1296 ( .A(n1457), .ZN(n1395) );
  NAND2_X1 U1297 ( .A1(n1402), .A2(n1404), .ZN(n768) );
  NOR2_X1 U1298 ( .A1(n1393), .A2(n610), .ZN(n1452) );
  AOI21_X2 U1304 ( .B1(n752), .B2(n735), .A(n1081), .ZN(n1116) );
  BUF_X4 U1305 ( .A(n968), .Z(n755) );
  NAND2_X2 U1307 ( .A1(n1028), .A2(n757), .ZN(n760) );
  NAND2_X2 U1308 ( .A1(n1629), .A2(n1464), .ZN(n1467) );
  BUF_X4 U1309 ( .A(n1153), .Z(n758) );
  NOR3_X2 U1310 ( .A1(n759), .A2(n1330), .A3(n1331), .ZN(\d[20] ) );
  NOR2_X2 U1311 ( .A1(n549), .A2(n712), .ZN(n759) );
  INV_X2 U1312 ( .A(n764), .ZN(n763) );
  NAND2_X1 U1315 ( .A1(n718), .A2(n1403), .ZN(n1333) );
  BUF_X4 U1317 ( .A(n945), .Z(n767) );
  OAI22_X2 U1319 ( .A1(n1489), .A2(n1625), .B1(n1491), .B2(n767), .ZN(n1494)
         );
  NAND2_X2 U1320 ( .A1(n873), .A2(n872), .ZN(n770) );
  NAND2_X1 U1322 ( .A1(n1545), .A2(n1495), .ZN(n1498) );
  AOI22_X2 U1326 ( .A1(n789), .A2(n1246), .B1(n1244), .B2(n1245), .ZN(n1283)
         );
  NAND3_X2 U1329 ( .A1(n905), .A2(n977), .A3(n976), .ZN(n793) );
  BUF_X4 U1331 ( .A(n1609), .Z(n798) );
  BUF_X4 U1336 ( .A(n820), .Z(n802) );
  NAND2_X1 U1337 ( .A1(n695), .A2(n820), .ZN(n1010) );
  NAND2_X1 U1338 ( .A1(n928), .A2(n820), .ZN(n935) );
  MUX2_X2 U1339 ( .A(n802), .B(n1376), .S(a[24]), .Z(n1371) );
  MUX2_X2 U1340 ( .A(n802), .B(n1376), .S(a[25]), .Z(n1377) );
  NAND2_X4 U1341 ( .A1(n1683), .A2(b[14]), .ZN(n820) );
  NAND2_X4 U1342 ( .A1(n687), .A2(n942), .ZN(n1033) );
  INV_X4 U1343 ( .A(n803), .ZN(n1118) );
  INV_X4 U1345 ( .A(n1118), .ZN(n804) );
  INV_X8 U1346 ( .A(n806), .ZN(n808) );
  NAND2_X2 U1347 ( .A1(n1263), .A2(n625), .ZN(n810) );
  NAND2_X2 U1348 ( .A1(n1054), .A2(n776), .ZN(n811) );
  NOR2_X2 U1350 ( .A1(n1066), .A2(n1065), .ZN(n814) );
  NAND2_X1 U1351 ( .A1(n505), .A2(n802), .ZN(n889) );
  NOR2_X4 U1352 ( .A1(n576), .A2(n1095), .ZN(n1100) );
  NAND2_X2 U1353 ( .A1(n1300), .A2(n1301), .ZN(n1334) );
  NAND2_X2 U1355 ( .A1(n831), .A2(n830), .ZN(n1262) );
  NAND2_X1 U1356 ( .A1(n257), .A2(n1412), .ZN(n830) );
  NAND2_X2 U1357 ( .A1(n282), .A2(n994), .ZN(n831) );
  NAND2_X1 U1358 ( .A1(n1047), .A2(n738), .ZN(n964) );
  NOR2_X4 U1359 ( .A1(n1038), .A2(n1039), .ZN(n1093) );
  NAND2_X2 U1360 ( .A1(n834), .A2(n833), .ZN(n1132) );
  NAND2_X2 U1361 ( .A1(n758), .A2(n1054), .ZN(n834) );
  BUF_X4 U1362 ( .A(n1710), .Z(n835) );
  BUF_X4 U1364 ( .A(n844), .Z(n837) );
  INV_X4 U1368 ( .A(n948), .ZN(n1263) );
  NAND2_X1 U1369 ( .A1(n947), .A2(n1412), .ZN(n1413) );
  NOR2_X1 U1372 ( .A1(n1454), .A2(n600), .ZN(n1455) );
  INV_X1 U1373 ( .A(n848), .ZN(n1014) );
  BUF_X4 U1375 ( .A(n97), .Z(n851) );
  AOI22_X2 U1380 ( .A1(n940), .A2(n546), .B1(n939), .B2(n550), .ZN(\d[19] ) );
  NOR2_X4 U1382 ( .A1(n1170), .A2(n1169), .ZN(n1175) );
  INV_X4 U1383 ( .A(n1467), .ZN(n869) );
  NAND2_X2 U1385 ( .A1(n949), .A2(n606), .ZN(n876) );
  NAND2_X2 U1388 ( .A1(n883), .A2(n882), .ZN(n881) );
  NAND2_X2 U1389 ( .A1(n802), .A2(n40), .ZN(n882) );
  NAND2_X2 U1390 ( .A1(n1376), .A2(n1160), .ZN(n883) );
  NOR2_X2 U1391 ( .A1(n885), .A2(n663), .ZN(n884) );
  NAND2_X2 U1393 ( .A1(n1470), .A2(n1471), .ZN(\d[13] ) );
  NAND2_X2 U1394 ( .A1(n890), .A2(n889), .ZN(n1156) );
  NAND2_X2 U1395 ( .A1(n1376), .A2(n625), .ZN(n890) );
  NAND2_X2 U1396 ( .A1(n1123), .A2(n1124), .ZN(n1150) );
  AOI22_X2 U1397 ( .A1(n1145), .A2(n1175), .B1(n1143), .B2(n1144), .ZN(n1182)
         );
  NOR2_X1 U1400 ( .A1(n558), .A2(n1420), .ZN(n1433) );
  NOR2_X1 U1401 ( .A1(n1261), .A2(n902), .ZN(n1260) );
  NAND2_X2 U1406 ( .A1(n917), .A2(n1219), .ZN(n940) );
  NAND2_X2 U1407 ( .A1(n920), .A2(n919), .ZN(n1299) );
  NAND2_X2 U1409 ( .A1(n925), .A2(n924), .ZN(n923) );
  NAND2_X2 U1410 ( .A1(n1614), .A2(n1400), .ZN(n1404) );
  BUF_X4 U1411 ( .A(n930), .Z(n929) );
  XNOR2_X1 U1412 ( .A(n929), .B(n1465), .ZN(n1466) );
  INV_X4 U1417 ( .A(n1286), .ZN(n945) );
  NAND2_X2 U1419 ( .A1(n1089), .A2(n1090), .ZN(n949) );
  INV_X2 U1420 ( .A(n1147), .ZN(n1300) );
  XOR2_X1 U1423 ( .A(n808), .B(a[20]), .Z(n1058) );
  XOR2_X1 U1424 ( .A(n808), .B(n1160), .Z(n1161) );
  INV_X8 U1427 ( .A(b[8]), .ZN(n1410) );
  XNOR2_X1 U1428 ( .A(n1209), .B(a[13]), .ZN(n1210) );
  XNOR2_X1 U1429 ( .A(n1209), .B(a[15]), .ZN(n969) );
  AND2_X4 U1430 ( .A1(n628), .A2(n1356), .ZN(n956) );
  INV_X2 U1431 ( .A(n1219), .ZN(n1497) );
  INV_X2 U1433 ( .A(n1089), .ZN(n1091) );
  NOR3_X1 U1434 ( .A1(n1232), .A2(n29), .A3(n1235), .ZN(n1233) );
  NAND2_X1 U1435 ( .A1(n1382), .A2(n45), .ZN(n1383) );
  INV_X1 U1436 ( .A(n1268), .ZN(n1266) );
  AOI21_X1 U1437 ( .B1(n1442), .B2(n1447), .A(n1430), .ZN(n1431) );
  AOI21_X1 U1438 ( .B1(n1434), .B2(n1436), .A(n1433), .ZN(n1421) );
  OAI21_X1 U1439 ( .B1(n1411), .B2(n1746), .A(a[8]), .ZN(n1415) );
  INV_X4 U1440 ( .A(b[11]), .ZN(n961) );
  INV_X4 U1441 ( .A(n961), .ZN(n1209) );
  INV_X8 U1442 ( .A(n618), .ZN(n1053) );
  INV_X8 U1443 ( .A(n961), .ZN(n968) );
  XNOR2_X2 U1444 ( .A(n989), .B(n1239), .ZN(n967) );
  NAND2_X2 U1445 ( .A1(n695), .A2(n808), .ZN(n971) );
  BUF_X4 U1446 ( .A(n1130), .Z(n1265) );
  INV_X8 U1447 ( .A(n806), .ZN(n989) );
  NAND2_X2 U1449 ( .A1(n970), .A2(n971), .ZN(n975) );
  BUF_X4 U1450 ( .A(a[16]), .Z(n1060) );
  BUF_X4 U1451 ( .A(n937), .Z(n1376) );
  INV_X4 U1452 ( .A(a[17]), .ZN(n1074) );
  NAND2_X2 U1453 ( .A1(a[12]), .A2(n805), .ZN(n988) );
  NAND2_X2 U1458 ( .A1(n998), .A2(n841), .ZN(n999) );
  NAND3_X2 U1459 ( .A1(n1017), .A2(n1016), .A3(n1015), .ZN(n1020) );
  NOR2_X2 U1460 ( .A1(n1023), .A2(n807), .ZN(n1024) );
  NOR2_X4 U1461 ( .A1(n1025), .A2(n1024), .ZN(n1095) );
  BUF_X4 U1463 ( .A(a[21]), .Z(n1160) );
  NAND2_X2 U1464 ( .A1(n40), .A2(n1509), .ZN(n1073) );
  NAND2_X2 U1465 ( .A1(n732), .A2(n1512), .ZN(n1061) );
  BUF_X4 U1466 ( .A(a[23]), .Z(n1164) );
  NAND2_X2 U1467 ( .A1(n1069), .A2(n1068), .ZN(n1070) );
  BUF_X4 U1469 ( .A(n1628), .Z(n1085) );
  INV_X2 U1473 ( .A(a[24]), .ZN(n1125) );
  XNOR2_X2 U1474 ( .A(n1209), .B(a[25]), .ZN(n1134) );
  NOR2_X4 U1476 ( .A1(n1137), .A2(n1138), .ZN(n1170) );
  NAND2_X2 U1477 ( .A1(n952), .A2(n460), .ZN(n1139) );
  NAND2_X2 U1478 ( .A1(n937), .A2(a[20]), .ZN(n1142) );
  MUX2_X2 U1480 ( .A(n758), .B(n20), .S(a[24]), .Z(n1154) );
  INV_X2 U1482 ( .A(n602), .ZN(n1159) );
  INV_X4 U1483 ( .A(n1175), .ZN(n1172) );
  OAI21_X2 U1485 ( .B1(n647), .B2(n794), .A(n493), .ZN(n1181) );
  NAND2_X2 U1486 ( .A1(n647), .A2(n794), .ZN(n1180) );
  INV_X4 U1487 ( .A(n1222), .ZN(n1216) );
  BUF_X4 U1488 ( .A(n1218), .Z(n1219) );
  BUF_X4 U1489 ( .A(n1234), .Z(n1228) );
  OAI21_X2 U1491 ( .B1(n461), .B2(n1260), .A(n1259), .ZN(n1436) );
  INV_X4 U1492 ( .A(n1269), .ZN(n1272) );
  NOR2_X2 U1493 ( .A1(n1274), .A2(n1273), .ZN(n1424) );
  INV_X4 U1495 ( .A(n1443), .ZN(n1441) );
  MUX2_X2 U1497 ( .A(n1303), .B(n1302), .S(a[25]), .Z(n1370) );
  NOR2_X1 U1498 ( .A1(n1305), .A2(n51), .ZN(n1307) );
  INV_X4 U1501 ( .A(n1323), .ZN(n1325) );
  AOI21_X2 U1502 ( .B1(n885), .B2(n663), .A(n1325), .ZN(n1327) );
  NOR2_X2 U1503 ( .A1(n1327), .A2(n1326), .ZN(n1331) );
  BUF_X4 U1507 ( .A(n1352), .Z(n1353) );
  NAND2_X2 U1510 ( .A1(n1375), .A2(n1374), .ZN(n1378) );
  INV_X2 U1511 ( .A(n1380), .ZN(n1381) );
  MUX2_X2 U1512 ( .A(n1383), .B(n1382), .S(n1381), .Z(n1388) );
  XNOR2_X2 U1515 ( .A(n1456), .B(n1455), .ZN(\d[9] ) );
  NAND2_X2 U1519 ( .A1(n1486), .A2(n1504), .ZN(n1488) );
  INV_X4 U1520 ( .A(n1488), .ZN(n1491) );
  NAND2_X2 U430 ( .A1(n901), .A2(n471), .ZN(n467) );
  INV_X4 U105 ( .A(n18), .ZN(n732) );
  NAND2_X4 U307 ( .A1(n875), .A2(n876), .ZN(n1088) );
  INV_X4 U175 ( .A(n443), .ZN(n177) );
  NOR2_X2 U309 ( .A1(n118), .A2(n689), .ZN(n1002) );
  INV_X4 U211 ( .A(n1237), .ZN(n47) );
  NAND2_X4 U934 ( .A1(n457), .A2(n454), .ZN(n1212) );
  NAND2_X2 U1194 ( .A1(n257), .A2(a[17]), .ZN(n1029) );
  NAND2_X2 U1131 ( .A1(n257), .A2(a[12]), .ZN(n580) );
  INV_X2 U906 ( .A(n428), .ZN(n427) );
  XNOR2_X2 U1425 ( .A(n805), .B(a[17]), .ZN(n1043) );
  INV_X4 U1010 ( .A(n1097), .ZN(n1094) );
  NOR2_X2 U1233 ( .A1(b[10]), .A2(n1053), .ZN(n1040) );
  INV_X4 U542 ( .A(n1108), .ZN(n692) );
  NAND2_X2 U253 ( .A1(n286), .A2(n1605), .ZN(n924) );
  INV_X4 U1260 ( .A(n1511), .ZN(n701) );
  NAND2_X2 U422 ( .A1(n230), .A2(n754), .ZN(n870) );
  INV_X4 U926 ( .A(n446), .ZN(n445) );
  NAND2_X2 U870 ( .A1(n987), .A2(n848), .ZN(n401) );
  NOR2_X4 U647 ( .A1(n1519), .A2(n848), .ZN(n850) );
  NAND2_X2 U152 ( .A1(n991), .A2(n807), .ZN(n992) );
  INV_X4 U440 ( .A(n937), .ZN(n350) );
  OAI21_X2 U133 ( .B1(n1151), .B2(n1150), .A(n644), .ZN(n920) );
  INV_X1 U1279 ( .A(n1156), .ZN(n717) );
  NOR2_X2 U1392 ( .A1(n1210), .A2(n887), .ZN(n1214) );
  NOR2_X2 U401 ( .A1(n119), .A2(n1209), .ZN(n118) );
  INV_X8 U941 ( .A(n799), .ZN(n460) );
  NAND2_X2 U848 ( .A1(n384), .A2(n383), .ZN(n1237) );
  NAND2_X2 U360 ( .A1(n601), .A2(n1632), .ZN(n95) );
  INV_X8 U1333 ( .A(n1053), .ZN(n799) );
  AOI21_X2 U1122 ( .B1(n57), .B2(n1746), .A(n573), .ZN(n572) );
  NAND2_X2 U606 ( .A1(n1192), .A2(n1655), .ZN(n200) );
  NAND2_X2 U866 ( .A1(n1505), .A2(n493), .ZN(n398) );
  NOR2_X4 U1133 ( .A1(n1215), .A2(n1214), .ZN(n1235) );
  INV_X4 U223 ( .A(n706), .ZN(n1127) );
  INV_X8 U1301 ( .A(n1065), .ZN(n757) );
  INV_X4 U466 ( .A(n817), .ZN(n137) );
  NAND2_X2 U171 ( .A1(n286), .A2(n1527), .ZN(n764) );
  NOR2_X2 U1500 ( .A1(n1540), .A2(n1321), .ZN(n1328) );
  INV_X4 U1306 ( .A(n1257), .ZN(n887) );
  INV_X2 U143 ( .A(a[20]), .ZN(n1140) );
  INV_X2 U1475 ( .A(n1134), .ZN(n1129) );
  INV_X2 U1295 ( .A(n894), .ZN(n1079) );
  INV_X2 U1494 ( .A(n1276), .ZN(n1277) );
  NOR2_X2 U29 ( .A1(n1133), .A2(n1132), .ZN(n1183) );
  NAND2_X2 U1415 ( .A1(n543), .A2(n1297), .ZN(n1495) );
  INV_X1 U1092 ( .A(n1354), .ZN(n665) );
  XNOR2_X1 U1514 ( .A(n1436), .B(n1437), .ZN(\d[6] ) );
  INV_X2 U58 ( .A(n1334), .ZN(n1321) );
  INV_X2 U186 ( .A(n1478), .ZN(n1479) );
  INV_X2 U130 ( .A(n1188), .ZN(n87) );
  INV_X2 U652 ( .A(n243), .ZN(n239) );
  INV_X2 U1105 ( .A(n1105), .ZN(n727) );
  NAND2_X2 U21 ( .A1(n1631), .A2(n727), .ZN(n1104) );
  BUF_X4 U187 ( .A(n1365), .Z(n159) );
  INV_X2 U89 ( .A(n159), .ZN(n1366) );
  INV_X4 U1115 ( .A(n560), .ZN(n559) );
  NAND2_X4 U47 ( .A1(n465), .A2(n464), .ZN(n1148) );
  INV_X4 U978 ( .A(n815), .ZN(n495) );
  NAND2_X2 U358 ( .A1(n1000), .A2(n999), .ZN(n1289) );
  NAND2_X2 U463 ( .A1(n1131), .A2(a[11]), .ZN(n228) );
  INV_X2 U1 ( .A(n124), .ZN(n1547) );
  INV_X4 U2 ( .A(n1052), .ZN(n1578) );
  INV_X4 U10 ( .A(n750), .ZN(n1606) );
  NAND2_X2 U25 ( .A1(n1270), .A2(n283), .ZN(n285) );
  NAND2_X1 U27 ( .A1(n1270), .A2(n1750), .ZN(n11) );
  NAND2_X1 U31 ( .A1(n55), .A2(n1703), .ZN(n79) );
  INV_X4 U32 ( .A(n704), .ZN(n1550) );
  INV_X2 U35 ( .A(n1520), .ZN(n746) );
  NAND2_X2 U39 ( .A1(n1550), .A2(n137), .ZN(n630) );
  INV_X1 U42 ( .A(n1019), .ZN(n1016) );
  NAND2_X2 U49 ( .A1(n55), .A2(n1529), .ZN(n180) );
  XOR2_X2 U51 ( .A(n808), .B(a[11]), .Z(n1203) );
  NAND2_X1 U53 ( .A1(n412), .A2(n822), .ZN(n145) );
  NAND2_X2 U59 ( .A1(n1243), .A2(n412), .ZN(n1251) );
  NAND2_X1 U60 ( .A1(n283), .A2(n412), .ZN(n1252) );
  NAND2_X1 U61 ( .A1(n412), .A2(n1750), .ZN(n1206) );
  NOR2_X4 U68 ( .A1(n1317), .A2(n89), .ZN(n1318) );
  INV_X4 U75 ( .A(n856), .ZN(n680) );
  NAND2_X4 U76 ( .A1(n84), .A2(n1140), .ZN(n855) );
  INV_X2 U84 ( .A(n600), .ZN(n1356) );
  NAND2_X2 U86 ( .A1(n1163), .A2(n1162), .ZN(n493) );
  NAND2_X2 U87 ( .A1(n523), .A2(n521), .ZN(n1097) );
  INV_X2 U88 ( .A(a[22]), .ZN(n1054) );
  INV_X2 U93 ( .A(n1348), .ZN(n1503) );
  INV_X2 U94 ( .A(n1285), .ZN(n1504) );
  NAND2_X2 U95 ( .A1(n447), .A2(n445), .ZN(n617) );
  INV_X2 U99 ( .A(n1230), .ZN(n1292) );
  NAND2_X2 U100 ( .A1(n88), .A2(n87), .ZN(n86) );
  INV_X2 U117 ( .A(n904), .ZN(n1588) );
  NAND2_X2 U120 ( .A1(n1563), .A2(n983), .ZN(n984) );
  NAND2_X2 U121 ( .A1(n653), .A2(n652), .ZN(n993) );
  INV_X4 U127 ( .A(n151), .ZN(n1508) );
  INV_X4 U137 ( .A(n1241), .ZN(n1509) );
  INV_X4 U139 ( .A(n1209), .ZN(n1510) );
  INV_X8 U144 ( .A(n618), .ZN(n1511) );
  INV_X4 U147 ( .A(n1060), .ZN(n1512) );
  NOR2_X4 U149 ( .A1(n1262), .A2(n9), .ZN(n1269) );
  NAND2_X1 U150 ( .A1(n756), .A2(n978), .ZN(n1515) );
  INV_X1 U158 ( .A(n756), .ZN(n1513) );
  AOI21_X2 U161 ( .B1(n947), .B2(a[12]), .A(n847), .ZN(n846) );
  NOR2_X1 U163 ( .A1(a[12]), .A2(n776), .ZN(n847) );
  XNOR2_X2 U182 ( .A(n1209), .B(n840), .ZN(n839) );
  INV_X2 U196 ( .A(n657), .ZN(n637) );
  AOI22_X1 U197 ( .A1(b[8]), .A2(n1012), .B1(n928), .B2(n1055), .ZN(n1517) );
  NAND2_X2 U199 ( .A1(n137), .A2(n1550), .ZN(n1518) );
  NAND2_X2 U203 ( .A1(n630), .A2(n156), .ZN(n1555) );
  NAND2_X2 U206 ( .A1(n102), .A2(n713), .ZN(n836) );
  NAND2_X2 U212 ( .A1(n321), .A2(n1662), .ZN(n296) );
  NAND2_X2 U214 ( .A1(n1213), .A2(n1212), .ZN(n1519) );
  NAND2_X2 U215 ( .A1(n1212), .A2(n1213), .ZN(n987) );
  INV_X2 U217 ( .A(n808), .ZN(n472) );
  AOI21_X2 U219 ( .B1(n307), .B2(n1289), .A(n1288), .ZN(n1520) );
  AOI22_X2 U226 ( .A1(n540), .A2(n724), .B1(n539), .B2(n723), .ZN(n1538) );
  NOR2_X1 U234 ( .A1(n1399), .A2(n97), .ZN(n1402) );
  NAND2_X2 U237 ( .A1(n1193), .A2(n50), .ZN(n1195) );
  NAND2_X2 U260 ( .A1(n504), .A2(n503), .ZN(n1165) );
  INV_X2 U265 ( .A(n986), .ZN(n578) );
  NOR3_X4 U266 ( .A1(n797), .A2(n1191), .A3(n1190), .ZN(n796) );
  NOR2_X4 U268 ( .A1(n367), .A2(n31), .ZN(n1191) );
  NAND2_X1 U271 ( .A1(n805), .A2(a[15]), .ZN(n1525) );
  NAND2_X1 U281 ( .A1(n1056), .A2(n1082), .ZN(n1083) );
  NOR2_X2 U282 ( .A1(n1364), .A2(n600), .ZN(n16) );
  NAND2_X1 U288 ( .A1(n1637), .A2(n1587), .ZN(n134) );
  INV_X1 U290 ( .A(n1403), .ZN(n1527) );
  NAND2_X2 U292 ( .A1(n991), .A2(n755), .ZN(n75) );
  NAND2_X1 U300 ( .A1(n1722), .A2(n1292), .ZN(n1394) );
  AND2_X2 U301 ( .A1(n1000), .A2(n999), .ZN(n1528) );
  INV_X2 U303 ( .A(n84), .ZN(n1529) );
  NAND2_X1 U304 ( .A1(n914), .A2(n1051), .ZN(n1114) );
  NAND2_X1 U314 ( .A1(n587), .A2(n722), .ZN(n326) );
  NAND2_X1 U316 ( .A1(n1531), .A2(n576), .ZN(n1532) );
  NAND2_X2 U318 ( .A1(n1530), .A2(n1095), .ZN(n1533) );
  NAND2_X2 U320 ( .A1(n1532), .A2(n1533), .ZN(n1034) );
  INV_X2 U321 ( .A(n576), .ZN(n1530) );
  INV_X1 U322 ( .A(n1095), .ZN(n1531) );
  INV_X2 U326 ( .A(n1034), .ZN(n149) );
  NAND2_X1 U328 ( .A1(n311), .A2(n1251), .ZN(n1536) );
  NAND2_X2 U330 ( .A1(n1534), .A2(n312), .ZN(n1537) );
  NAND2_X2 U331 ( .A1(n1536), .A2(n1537), .ZN(n168) );
  INV_X2 U343 ( .A(n311), .ZN(n1534) );
  NAND2_X1 U353 ( .A1(n357), .A2(n654), .ZN(n356) );
  NAND2_X1 U355 ( .A1(n155), .A2(n327), .ZN(n1554) );
  INV_X2 U362 ( .A(n70), .ZN(n69) );
  NAND2_X1 U365 ( .A1(n741), .A2(n1227), .ZN(n669) );
  NAND2_X2 U366 ( .A1(n695), .A2(n84), .ZN(n997) );
  NAND3_X1 U397 ( .A1(n1401), .A2(n1659), .A3(n1344), .ZN(n1345) );
  INV_X4 U398 ( .A(n1186), .ZN(n157) );
  NAND2_X2 U421 ( .A1(n40), .A2(n591), .ZN(n353) );
  INV_X1 U423 ( .A(n631), .ZN(n1545) );
  INV_X4 U426 ( .A(n407), .ZN(n631) );
  INV_X1 U432 ( .A(n149), .ZN(n1620) );
  NAND2_X1 U434 ( .A1(n1167), .A2(n1083), .ZN(n587) );
  INV_X4 U438 ( .A(n1403), .ZN(n1472) );
  NAND2_X1 U446 ( .A1(n675), .A2(n704), .ZN(n1552) );
  NAND2_X2 U450 ( .A1(n1551), .A2(n1550), .ZN(n1553) );
  NAND2_X2 U452 ( .A1(n1552), .A2(n1553), .ZN(n1032) );
  INV_X1 U453 ( .A(n675), .ZN(n1551) );
  NAND2_X1 U454 ( .A1(n558), .A2(n1420), .ZN(n1434) );
  NAND2_X2 U458 ( .A1(n155), .A2(n327), .ZN(n300) );
  NAND2_X1 U460 ( .A1(n948), .A2(a[24]), .ZN(n1068) );
  NAND2_X1 U461 ( .A1(n179), .A2(a[13]), .ZN(n996) );
  NAND2_X4 U465 ( .A1(n1261), .A2(n902), .ZN(n1259) );
  NAND2_X4 U468 ( .A1(n617), .A2(n616), .ZN(n605) );
  INV_X1 U472 ( .A(n1086), .ZN(n1614) );
  INV_X4 U477 ( .A(n989), .ZN(n689) );
  NAND2_X1 U482 ( .A1(n625), .A2(n160), .ZN(n503) );
  INV_X2 U483 ( .A(n468), .ZN(n901) );
  NAND2_X1 U485 ( .A1(n947), .A2(n1239), .ZN(n420) );
  NOR2_X1 U503 ( .A1(n1393), .A2(n1392), .ZN(n1637) );
  INV_X4 U506 ( .A(n1001), .ZN(n1239) );
  NAND2_X2 U510 ( .A1(n874), .A2(n1102), .ZN(n1580) );
  AOI21_X2 U516 ( .B1(n1079), .B2(n1080), .A(n1078), .ZN(n1102) );
  INV_X4 U517 ( .A(n174), .ZN(n173) );
  NAND2_X2 U527 ( .A1(n962), .A2(n1053), .ZN(n179) );
  NAND2_X2 U529 ( .A1(n900), .A2(n899), .ZN(n115) );
  NAND2_X2 U532 ( .A1(n1075), .A2(n757), .ZN(n900) );
  NAND3_X2 U535 ( .A1(n63), .A2(n1042), .A3(n1559), .ZN(n1098) );
  NAND2_X1 U538 ( .A1(n808), .A2(a[19]), .ZN(n1568) );
  NAND3_X2 U541 ( .A1(n116), .A2(n548), .A3(n175), .ZN(n1602) );
  INV_X4 U544 ( .A(n1560), .ZN(n877) );
  NAND2_X2 U549 ( .A1(n707), .A2(n136), .ZN(n1560) );
  NAND2_X2 U555 ( .A1(n704), .A2(n817), .ZN(n156) );
  NAND2_X2 U557 ( .A1(n1127), .A2(n1126), .ZN(n518) );
  INV_X4 U558 ( .A(n1022), .ZN(n1569) );
  NOR2_X4 U560 ( .A1(n1510), .A2(n1561), .ZN(n1131) );
  NAND2_X2 U561 ( .A1(b[12]), .A2(n1683), .ZN(n1561) );
  NAND2_X2 U567 ( .A1(n700), .A2(n1562), .ZN(n1636) );
  NAND2_X2 U569 ( .A1(n1223), .A2(n1237), .ZN(n1562) );
  NAND2_X2 U570 ( .A1(n900), .A2(n899), .ZN(n622) );
  NAND2_X2 U577 ( .A1(n937), .A2(a[11]), .ZN(n792) );
  INV_X2 U578 ( .A(n1633), .ZN(n193) );
  NAND2_X2 U584 ( .A1(n1570), .A2(n1571), .ZN(n117) );
  NOR2_X2 U585 ( .A1(n117), .A2(n1202), .ZN(n1288) );
  AOI22_X2 U601 ( .A1(n836), .A2(n640), .B1(n877), .B2(n1588), .ZN(n817) );
  NAND3_X2 U603 ( .A1(n1345), .A2(n1564), .A3(n1347), .ZN(n152) );
  AOI21_X2 U615 ( .B1(n488), .B2(n269), .A(n487), .ZN(n765) );
  INV_X2 U616 ( .A(n697), .ZN(n1593) );
  NAND2_X2 U617 ( .A1(n489), .A2(n695), .ZN(n697) );
  NAND2_X1 U619 ( .A1(a[13]), .A2(n1511), .ZN(n696) );
  NAND2_X2 U620 ( .A1(n775), .A2(n1218), .ZN(n719) );
  NAND2_X2 U628 ( .A1(n1368), .A2(n1367), .ZN(n1218) );
  NAND2_X2 U634 ( .A1(n273), .A2(a[18]), .ZN(n1563) );
  NAND2_X2 U635 ( .A1(n302), .A2(n677), .ZN(n679) );
  NAND2_X2 U636 ( .A1(n303), .A2(n305), .ZN(n302) );
  NAND2_X2 U644 ( .A1(n1481), .A2(n1625), .ZN(n1482) );
  NAND2_X2 U646 ( .A1(n292), .A2(n291), .ZN(n129) );
  NAND2_X2 U648 ( .A1(n955), .A2(n954), .ZN(n639) );
  NAND2_X2 U654 ( .A1(n963), .A2(n964), .ZN(n955) );
  NAND2_X2 U659 ( .A1(n400), .A2(n721), .ZN(n731) );
  NAND2_X2 U665 ( .A1(n101), .A2(n100), .ZN(n1643) );
  NAND2_X2 U666 ( .A1(n98), .A2(n102), .ZN(n101) );
  AND2_X2 U678 ( .A1(n1348), .A2(n1349), .ZN(n932) );
  NOR2_X2 U679 ( .A1(n1480), .A2(n782), .ZN(n781) );
  INV_X4 U685 ( .A(n1401), .ZN(n1480) );
  NOR2_X4 U688 ( .A1(n804), .A2(n868), .ZN(n1401) );
  AOI22_X2 U693 ( .A1(n229), .A2(n228), .B1(n226), .B2(n227), .ZN(n1632) );
  NAND2_X4 U694 ( .A1(n1153), .A2(n978), .ZN(n227) );
  INV_X2 U695 ( .A(n1184), .ZN(n773) );
  NAND2_X2 U699 ( .A1(n634), .A2(n633), .ZN(n1184) );
  INV_X2 U705 ( .A(n501), .ZN(n499) );
  NAND2_X2 U713 ( .A1(n710), .A2(n711), .ZN(n501) );
  XNOR2_X2 U716 ( .A(n1565), .B(n1359), .ZN(\d[10] ) );
  AOI22_X2 U721 ( .A1(n1566), .A2(n44), .B1(n322), .B2(n296), .ZN(n294) );
  NAND2_X2 U723 ( .A1(n1663), .A2(n1600), .ZN(n1566) );
  NAND2_X2 U727 ( .A1(n1567), .A2(n808), .ZN(n974) );
  NAND2_X2 U731 ( .A1(n468), .A2(n991), .ZN(n1567) );
  NAND2_X2 U737 ( .A1(n691), .A2(n1568), .ZN(n1066) );
  NAND2_X2 U739 ( .A1(n1569), .A2(n1001), .ZN(n615) );
  NAND2_X2 U741 ( .A1(n227), .A2(n226), .ZN(n1570) );
  NAND2_X2 U742 ( .A1(n228), .A2(n229), .ZN(n1571) );
  NAND2_X2 U745 ( .A1(n1158), .A2(n655), .ZN(n1572) );
  NOR2_X2 U751 ( .A1(n1660), .A2(n663), .ZN(n299) );
  NAND2_X2 U752 ( .A1(n1574), .A2(n1573), .ZN(n1155) );
  NAND2_X2 U753 ( .A1(n52), .A2(a[25]), .ZN(n1573) );
  NAND2_X2 U754 ( .A1(n1152), .A2(n952), .ZN(n1574) );
  NOR2_X1 U758 ( .A1(n602), .A2(n1384), .ZN(n1600) );
  AOI22_X2 U760 ( .A1(n1001), .A2(n591), .B1(n257), .B2(n1239), .ZN(n402) );
  NAND2_X2 U762 ( .A1(a[15]), .A2(n1053), .ZN(n652) );
  NAND2_X2 U770 ( .A1(n1349), .A2(n1337), .ZN(n602) );
  INV_X2 U772 ( .A(n1387), .ZN(n184) );
  NAND2_X2 U775 ( .A1(n185), .A2(n1337), .ZN(n1387) );
  NAND2_X2 U786 ( .A1(n893), .A2(n1657), .ZN(n895) );
  NAND3_X2 U798 ( .A1(n1612), .A2(n236), .A3(n235), .ZN(n234) );
  NAND2_X2 U802 ( .A1(n1577), .A2(n1394), .ZN(n316) );
  NAND3_X2 U810 ( .A1(n1721), .A2(n89), .A3(n628), .ZN(n103) );
  AOI22_X2 U814 ( .A1(n1107), .A2(n1104), .B1(n1684), .B2(n1105), .ZN(n750) );
  NAND2_X2 U818 ( .A1(n1621), .A2(n512), .ZN(n1457) );
  AOI21_X2 U821 ( .B1(n176), .B2(n1020), .A(n442), .ZN(n1627) );
  NOR2_X2 U830 ( .A1(n1276), .A2(n1275), .ZN(n1425) );
  AOI22_X2 U835 ( .A1(n1101), .A2(n749), .B1(n754), .B2(n1108), .ZN(n1631) );
  NAND2_X2 U844 ( .A1(n1259), .A2(n248), .ZN(n166) );
  INV_X4 U845 ( .A(n655), .ZN(n826) );
  NOR2_X2 U846 ( .A1(n1720), .A2(n1622), .ZN(n1630) );
  NAND2_X2 U857 ( .A1(n1578), .A2(n335), .ZN(n547) );
  NOR2_X4 U858 ( .A1(n1111), .A2(n1109), .ZN(n1052) );
  NAND2_X2 U862 ( .A1(n1613), .A2(n1209), .ZN(n65) );
  AOI21_X2 U867 ( .B1(n1046), .B2(b[8]), .A(n1045), .ZN(n1607) );
  INV_X2 U878 ( .A(n766), .ZN(n1579) );
  NAND2_X4 U880 ( .A1(n1511), .A2(n1410), .ZN(n1241) );
  OAI21_X2 U885 ( .B1(n1624), .B2(n1655), .A(n202), .ZN(n201) );
  NAND2_X2 U895 ( .A1(n481), .A2(n480), .ZN(n1624) );
  OAI21_X1 U896 ( .B1(n993), .B2(n1410), .A(n1508), .ZN(n741) );
  NAND2_X4 U897 ( .A1(n1511), .A2(n1410), .ZN(n1609) );
  NOR2_X4 U900 ( .A1(n1609), .A2(n1239), .ZN(n151) );
  NAND3_X2 U909 ( .A1(n816), .A2(n1732), .A3(n1251), .ZN(n1597) );
  NAND2_X2 U912 ( .A1(n495), .A2(n507), .ZN(n816) );
  NAND2_X2 U914 ( .A1(n796), .A2(n1624), .ZN(n583) );
  NAND2_X2 U915 ( .A1(n754), .A2(n1108), .ZN(n1603) );
  NAND2_X2 U938 ( .A1(n1100), .A2(n1710), .ZN(n1585) );
  BUF_X4 U954 ( .A(n869), .Z(n1586) );
  NOR2_X2 U965 ( .A1(n1720), .A2(n1622), .ZN(n1379) );
  NAND2_X2 U976 ( .A1(n1509), .A2(n1047), .ZN(n454) );
  AOI22_X2 U980 ( .A1(b[8]), .A2(n824), .B1(n1509), .B2(n822), .ZN(n1096) );
  NAND2_X4 U986 ( .A1(n620), .A2(n619), .ZN(n1257) );
  NAND2_X1 U991 ( .A1(n551), .A2(n1394), .ZN(n1587) );
  NOR2_X1 U994 ( .A1(a[17]), .A2(n1410), .ZN(n22) );
  NOR3_X4 U998 ( .A1(n1286), .A2(n1285), .A3(n1403), .ZN(n89) );
  NAND2_X2 U1004 ( .A1(n757), .A2(n967), .ZN(n136) );
  NAND2_X2 U1005 ( .A1(n845), .A2(a[17]), .ZN(n1006) );
  NOR2_X2 U1008 ( .A1(n968), .A2(b[12]), .ZN(n109) );
  NAND2_X2 U1011 ( .A1(n294), .A2(n295), .ZN(n293) );
  NAND2_X2 U1025 ( .A1(n1340), .A2(n1589), .ZN(n139) );
  INV_X2 U1028 ( .A(n1332), .ZN(n1591) );
  NAND2_X2 U1031 ( .A1(n841), .A2(n839), .ZN(n351) );
  NOR2_X2 U1035 ( .A1(n1594), .A2(n1593), .ZN(n222) );
  NAND2_X2 U1038 ( .A1(n696), .A2(b[8]), .ZN(n1594) );
  NAND2_X2 U1043 ( .A1(n1595), .A2(n1052), .ZN(n745) );
  AOI22_X2 U1045 ( .A1(n686), .A2(n687), .B1(n914), .B2(n1051), .ZN(n335) );
  INV_X4 U1053 ( .A(n738), .ZN(n995) );
  XNOR2_X2 U1055 ( .A(n756), .B(n1596), .ZN(n998) );
  INV_X2 U1058 ( .A(n1239), .ZN(n1596) );
  NAND3_X2 U1076 ( .A1(n1597), .A2(n310), .A3(n308), .ZN(n343) );
  NAND2_X2 U1084 ( .A1(n881), .A2(n655), .ZN(n533) );
  AND2_X2 U1085 ( .A1(n989), .A2(a[10]), .ZN(n450) );
  OAI21_X2 U1102 ( .B1(n224), .B2(n807), .A(n1601), .ZN(n1227) );
  XNOR2_X2 U1127 ( .A(n1053), .B(n801), .ZN(n824) );
  NAND2_X2 U1129 ( .A1(n1638), .A2(n1602), .ZN(\d[17] ) );
  NAND2_X2 U1134 ( .A1(n1604), .A2(n1603), .ZN(n1647) );
  NAND2_X2 U1135 ( .A1(n749), .A2(n1101), .ZN(n1604) );
  INV_X1 U1138 ( .A(n138), .ZN(n1362) );
  INV_X4 U1139 ( .A(n1189), .ZN(n368) );
  INV_X1 U1140 ( .A(n1294), .ZN(n705) );
  AND2_X2 U1141 ( .A1(n597), .A2(n411), .ZN(n35) );
  NAND2_X1 U1149 ( .A1(n1487), .A2(n1459), .ZN(n1463) );
  NAND2_X1 U1156 ( .A1(n1060), .A2(n1131), .ZN(n1042) );
  NAND2_X1 U1157 ( .A1(n1472), .A2(n97), .ZN(n1605) );
  NAND2_X2 U1165 ( .A1(n97), .A2(n1472), .ZN(n59) );
  NAND2_X1 U1172 ( .A1(n1140), .A2(n394), .ZN(n1080) );
  NAND2_X4 U1173 ( .A1(n1055), .A2(n1512), .ZN(n905) );
  NAND2_X1 U1174 ( .A1(n1389), .A2(n1344), .ZN(n1347) );
  INV_X2 U1179 ( .A(n1389), .ZN(n1342) );
  XNOR2_X2 U1181 ( .A(n288), .B(n1606), .ZN(n1475) );
  NAND2_X4 U1183 ( .A1(n458), .A2(b[8]), .ZN(n457) );
  NAND2_X1 U1193 ( .A1(n845), .A2(a[10]), .ZN(n10) );
  NAND2_X1 U1203 ( .A1(n845), .A2(n1164), .ZN(n78) );
  NAND2_X2 U1215 ( .A1(n951), .A2(n352), .ZN(n1608) );
  NAND2_X2 U1219 ( .A1(n352), .A2(n951), .ZN(n531) );
  NAND2_X1 U1220 ( .A1(n640), .A2(n836), .ZN(n207) );
  INV_X2 U1224 ( .A(n850), .ZN(n236) );
  INV_X2 U1235 ( .A(n1309), .ZN(n1310) );
  INV_X4 U1238 ( .A(n1086), .ZN(n718) );
  NAND2_X1 U1240 ( .A1(n623), .A2(n685), .ZN(n418) );
  NOR2_X2 U1245 ( .A1(n835), .A2(n30), .ZN(n436) );
  NAND2_X2 U1247 ( .A1(n178), .A2(n177), .ZN(n1615) );
  NAND2_X2 U1249 ( .A1(n178), .A2(n177), .ZN(n66) );
  NOR2_X4 U1252 ( .A1(n626), .A2(n1390), .ZN(n1616) );
  NOR2_X2 U1254 ( .A1(n626), .A2(n1390), .ZN(n1363) );
  INV_X2 U1256 ( .A(n1117), .ZN(n868) );
  NAND2_X2 U1270 ( .A1(n1284), .A2(n1418), .ZN(n1617) );
  NAND2_X1 U1283 ( .A1(n302), .A2(n677), .ZN(n1619) );
  INV_X2 U1287 ( .A(n639), .ZN(n98) );
  NAND3_X2 U1293 ( .A1(n399), .A2(n795), .A3(n398), .ZN(n480) );
  INV_X4 U1294 ( .A(n1107), .ZN(n435) );
  NAND2_X2 U1299 ( .A1(n66), .A2(n656), .ZN(n1621) );
  NAND2_X2 U1300 ( .A1(n1615), .A2(n656), .ZN(n1352) );
  NOR2_X2 U1302 ( .A1(n1099), .A2(n1098), .ZN(n749) );
  NAND2_X2 U1303 ( .A1(n17), .A2(n16), .ZN(n1622) );
  AND2_X4 U1316 ( .A1(n986), .A2(n211), .ZN(n1623) );
  NOR2_X4 U1321 ( .A1(n930), .A2(n1464), .ZN(n1286) );
  NOR2_X1 U1323 ( .A1(n37), .A2(n1616), .ZN(n332) );
  NAND2_X4 U1324 ( .A1(n278), .A2(n277), .ZN(n1107) );
  AOI21_X1 U1330 ( .B1(n1130), .B2(a[18]), .A(n808), .ZN(n1064) );
  NOR2_X2 U1334 ( .A1(n147), .A2(n1398), .ZN(n1625) );
  NOR2_X2 U1335 ( .A1(n1398), .A2(n147), .ZN(n1626) );
  NOR2_X2 U1354 ( .A1(n147), .A2(n1398), .ZN(n1490) );
  NAND2_X2 U1363 ( .A1(n1337), .A2(n1349), .ZN(n1385) );
  XNOR2_X2 U1365 ( .A(n1304), .B(n1373), .ZN(n1382) );
  INV_X4 U1370 ( .A(n1490), .ZN(n552) );
  NAND2_X1 U1374 ( .A1(n77), .A2(n1032), .ZN(n153) );
  NOR2_X1 U1376 ( .A1(n77), .A2(n1032), .ZN(n1031) );
  AOI21_X2 U1379 ( .B1(n874), .B2(n1102), .A(n766), .ZN(n1628) );
  NAND2_X4 U1381 ( .A1(n1199), .A2(n1198), .ZN(n1390) );
  NAND2_X2 U1384 ( .A1(n356), .A2(n677), .ZN(n1199) );
  NAND2_X1 U1399 ( .A1(n1018), .A2(n1643), .ZN(n515) );
  NOR3_X2 U1402 ( .A1(n364), .A2(n363), .A3(n368), .ZN(n1190) );
  NAND3_X2 U1408 ( .A1(n168), .A2(n1259), .A3(n248), .ZN(n167) );
  NAND2_X2 U1413 ( .A1(n679), .A2(n678), .ZN(n146) );
  NAND3_X2 U1414 ( .A1(n301), .A2(n303), .A3(n305), .ZN(n678) );
  NAND2_X2 U1432 ( .A1(n1635), .A2(n621), .ZN(n569) );
  NAND2_X2 U1454 ( .A1(n538), .A2(n1636), .ZN(n537) );
  NAND2_X2 U1462 ( .A1(n712), .A2(n1391), .ZN(n1638) );
  NAND2_X2 U1468 ( .A1(n1639), .A2(n256), .ZN(n556) );
  NOR2_X2 U1471 ( .A1(n819), .A2(n818), .ZN(n514) );
  NAND2_X2 U1479 ( .A1(n1640), .A2(n724), .ZN(n704) );
  NAND3_X2 U1496 ( .A1(n1641), .A2(n915), .A3(n313), .ZN(n248) );
  INV_X2 U1508 ( .A(n1296), .ZN(n1297) );
  NAND2_X1 U1509 ( .A1(n551), .A2(n1220), .ZN(n597) );
  INV_X2 U1516 ( .A(n741), .ZN(n667) );
  NAND2_X1 U1521 ( .A1(n389), .A2(n256), .ZN(n1644) );
  NAND2_X2 U1522 ( .A1(n256), .A2(n389), .ZN(n255) );
  NOR2_X2 U1524 ( .A1(n135), .A2(n97), .ZN(n1645) );
  NOR2_X2 U1525 ( .A1(n135), .A2(n97), .ZN(n1343) );
  NOR3_X1 U1526 ( .A1(n1644), .A2(n514), .A3(n254), .ZN(n1646) );
  NAND2_X2 U1528 ( .A1(n524), .A2(n1510), .ZN(n523) );
  BUF_X4 U1530 ( .A(n1197), .Z(n1649) );
  NAND2_X2 U1531 ( .A1(n1651), .A2(n1650), .ZN(n950) );
  INV_X2 U1532 ( .A(n1056), .ZN(n1650) );
  INV_X2 U1533 ( .A(n1082), .ZN(n1651) );
  NAND2_X2 U1535 ( .A1(n843), .A2(n1089), .ZN(n304) );
  INV_X4 U1537 ( .A(n1653), .ZN(n584) );
  NOR2_X2 U1538 ( .A1(n796), .A2(n1192), .ZN(n1653) );
  NAND2_X2 U1539 ( .A1(n1654), .A2(n362), .ZN(n797) );
  NAND2_X2 U1540 ( .A1(n361), .A2(n31), .ZN(n1654) );
  INV_X4 U1541 ( .A(n1474), .ZN(n288) );
  NAND2_X2 U1542 ( .A1(n400), .A2(n721), .ZN(n1474) );
  BUF_X4 U1543 ( .A(n364), .Z(n1655) );
  NOR2_X2 U1544 ( .A1(n1130), .A2(a[8]), .ZN(n91) );
  NAND3_X2 U1545 ( .A1(n25), .A2(n809), .A3(n941), .ZN(n939) );
  NAND2_X4 U1547 ( .A1(n1257), .A2(n755), .ZN(n394) );
  NAND2_X2 U1548 ( .A1(n1176), .A2(n676), .ZN(n866) );
  NAND2_X2 U1549 ( .A1(n778), .A2(n1656), .ZN(n1109) );
  NAND2_X1 U1550 ( .A1(n1270), .A2(n928), .ZN(n1656) );
  OR2_X2 U1551 ( .A1(n76), .A2(n75), .ZN(n1657) );
  INV_X1 U1552 ( .A(n1586), .ZN(n733) );
  NAND2_X4 U1553 ( .A1(n285), .A2(n83), .ZN(n1443) );
  INV_X2 U1554 ( .A(n1646), .ZN(n909) );
  INV_X4 U1555 ( .A(n359), .ZN(n17) );
  NOR2_X4 U1557 ( .A1(n1324), .A2(n1365), .ZN(n2) );
  NAND2_X2 U813 ( .A1(n1474), .A2(n750), .ZN(n1473) );
  INV_X1 U982 ( .A(n1257), .ZN(n76) );
  INV_X2 U785 ( .A(n895), .ZN(n853) );
  INV_X4 U1289 ( .A(b[10]), .ZN(n965) );
  INV_X8 U1403 ( .A(n903), .ZN(n937) );
  NOR2_X4 U310 ( .A1(b[14]), .A2(n1683), .ZN(n903) );
  NAND2_X2 U860 ( .A1(n1247), .A2(n1522), .ZN(n612) );
  INV_X4 U1236 ( .A(n1507), .ZN(n1612) );
  INV_X2 U755 ( .A(n1251), .ZN(n312) );
  AOI21_X2 U134 ( .B1(n746), .B2(n389), .A(n388), .ZN(n387) );
  NAND2_X2 U241 ( .A1(n312), .A2(n1247), .ZN(n310) );
  NAND2_X4 U939 ( .A1(n684), .A2(n683), .ZN(n458) );
  NAND2_X2 U1241 ( .A1(n751), .A2(n1511), .ZN(n683) );
  NAND2_X2 U1171 ( .A1(n1140), .A2(n820), .ZN(n1141) );
  INV_X4 U399 ( .A(n621), .ZN(n568) );
  INV_X4 U997 ( .A(n1100), .ZN(n1108) );
  INV_X4 U104 ( .A(n1179), .ZN(n1505) );
  INV_X4 U1029 ( .A(n536), .ZN(n535) );
  NAND2_X2 U269 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NAND2_X2 U1150 ( .A1(n780), .A2(n1146), .ZN(n592) );
  NOR2_X2 U364 ( .A1(n1009), .A2(n1008), .ZN(n540) );
  NOR2_X2 U136 ( .A1(n1480), .A2(n768), .ZN(n832) );
  NAND2_X4 U17 ( .A1(n86), .A2(n85), .ZN(n1197) );
  NAND2_X2 U373 ( .A1(n65), .A2(a[17]), .ZN(n938) );
  NAND2_X4 U1523 ( .A1(n1209), .A2(n965), .ZN(n459) );
  NAND2_X2 U1073 ( .A1(n625), .A2(n20), .ZN(n833) );
  INV_X1 U956 ( .A(n1183), .ZN(n648) );
  NAND2_X4 U960 ( .A1(n534), .A2(n533), .ZN(n780) );
  NAND2_X2 U148 ( .A1(n1115), .A2(n835), .ZN(n438) );
  INV_X2 U16 ( .A(n1094), .ZN(n872) );
  BUF_X4 U1151 ( .A(n1131), .Z(n20) );
  NAND2_X2 U1457 ( .A1(n997), .A2(n996), .ZN(n1000) );
  NAND2_X2 U374 ( .A1(a[10]), .A2(n65), .ZN(n1205) );
  INV_X2 U183 ( .A(n884), .ZN(n1329) );
  INV_X2 U254 ( .A(n1165), .ZN(n396) );
  NAND2_X2 U342 ( .A1(n84), .A2(n505), .ZN(n504) );
  INV_X2 U489 ( .A(n795), .ZN(n395) );
  NAND2_X2 U519 ( .A1(n40), .A2(n1511), .ZN(n1558) );
  INV_X2 U1024 ( .A(n780), .ZN(n532) );
  NAND2_X4 U1026 ( .A1(n826), .A2(n737), .ZN(n534) );
  AOI21_X2 U167 ( .B1(n1167), .B2(n1083), .A(n854), .ZN(n375) );
  OAI22_X2 U1422 ( .A1(n1626), .A2(n1469), .B1(n1586), .B2(n730), .ZN(n1470)
         );
  NAND2_X2 U1213 ( .A1(a[24]), .A2(n845), .ZN(n214) );
  INV_X1 U533 ( .A(n369), .ZN(n1158) );
  NAND2_X2 U1239 ( .A1(n1407), .A2(n1480), .ZN(n1409) );
  NOR3_X2 U687 ( .A1(n262), .A2(n1404), .A3(n1730), .ZN(n1407) );
  INV_X2 U82 ( .A(n914), .ZN(n686) );
  INV_X4 U118 ( .A(n849), .ZN(n1507) );
  INV_X2 U656 ( .A(n1115), .ZN(n245) );
  NOR2_X2 U868 ( .A1(n1748), .A2(n493), .ZN(n753) );
  NAND2_X2 U777 ( .A1(a[20]), .A2(n336), .ZN(n674) );
  NAND2_X2 U547 ( .A1(n1142), .A2(n1141), .ZN(n1174) );
  NAND2_X2 U129 ( .A1(n823), .A2(n821), .ZN(n1169) );
  NAND2_X2 U1405 ( .A1(n1255), .A2(n1256), .ZN(n915) );
  INV_X2 U520 ( .A(n1116), .ZN(n268) );
  INV_X2 U780 ( .A(n671), .ZN(n337) );
  INV_X2 U40 ( .A(n1436), .ZN(n1280) );
  INV_X1 U1090 ( .A(n1449), .ZN(n1442) );
  INV_X2 U1470 ( .A(n514), .ZN(n1639) );
  NOR2_X1 U85 ( .A1(n1498), .A2(n1497), .ZN(n550) );
  AND2_X1 U1101 ( .A1(n25), .A2(n1498), .ZN(n546) );
  INV_X2 U315 ( .A(n933), .ZN(n1350) );
  NOR2_X2 U674 ( .A1(n615), .A2(n253), .ZN(n1025) );
  NAND2_X2 U1034 ( .A1(n591), .A2(n1125), .ZN(n1126) );
  NOR2_X2 U5 ( .A1(n222), .A2(n815), .ZN(n311) );
  NOR2_X2 U1481 ( .A1(n1155), .A2(n1154), .ZN(n1373) );
  NOR2_X1 U966 ( .A1(n1447), .A2(n1424), .ZN(n486) );
  NOR2_X2 U4 ( .A1(n1494), .A2(n1493), .ZN(\d[14] ) );
  NAND2_X2 U13 ( .A1(n537), .A2(n535), .ZN(n1393) );
  NAND2_X4 U14 ( .A1(n1128), .A2(n1129), .ZN(n369) );
  OR2_X2 U18 ( .A1(n1385), .A2(n1386), .ZN(n1660) );
  AND3_X1 U22 ( .A1(n429), .A2(n36), .A3(n1159), .ZN(n1661) );
  AND3_X1 U23 ( .A1(n1495), .A2(n1336), .A3(n1334), .ZN(n1662) );
  INV_X2 U24 ( .A(n624), .ZN(n973) );
  INV_X4 U26 ( .A(n448), .ZN(n447) );
  NAND2_X4 U28 ( .A1(n968), .A2(b[12]), .ZN(n107) );
  NAND2_X4 U30 ( .A1(n500), .A2(n498), .ZN(n502) );
  NAND2_X4 U38 ( .A1(n703), .A2(n1558), .ZN(n1046) );
  INV_X8 U41 ( .A(n107), .ZN(n1130) );
  INV_X4 U46 ( .A(n343), .ZN(n342) );
  NAND2_X2 U52 ( .A1(n992), .A2(n93), .ZN(n229) );
  INV_X2 U67 ( .A(n1130), .ZN(n93) );
  INV_X4 U69 ( .A(n663), .ZN(n1663) );
  NAND2_X2 U73 ( .A1(n1010), .A2(n1011), .ZN(n943) );
  NOR2_X1 U77 ( .A1(n763), .A2(n851), .ZN(n1477) );
  INV_X2 U78 ( .A(n851), .ZN(n1486) );
  AND2_X1 U79 ( .A1(n1348), .A2(n1645), .ZN(n1659) );
  AND2_X1 U80 ( .A1(n1645), .A2(n1117), .ZN(n1669) );
  INV_X1 U81 ( .A(n1477), .ZN(n782) );
  AND2_X1 U83 ( .A1(n605), .A2(n1283), .ZN(n1502) );
  INV_X2 U96 ( .A(n566), .ZN(n1444) );
  NAND2_X2 U98 ( .A1(n1443), .A2(n566), .ZN(n1447) );
  NOR2_X2 U103 ( .A1(n566), .A2(n1443), .ZN(n1430) );
  NAND2_X2 U107 ( .A1(n734), .A2(n1645), .ZN(n1664) );
  NAND2_X1 U112 ( .A1(n1122), .A2(n757), .ZN(n1123) );
  NAND2_X1 U113 ( .A1(n1161), .A2(n757), .ZN(n1162) );
  NAND2_X1 U114 ( .A1(n1040), .A2(n928), .ZN(n522) );
  INV_X1 U123 ( .A(n1054), .ZN(n625) );
  NAND2_X1 U124 ( .A1(n591), .A2(n1512), .ZN(n828) );
  OR2_X1 U131 ( .A1(n466), .A2(n737), .ZN(n32) );
  XOR2_X1 U145 ( .A(n780), .B(n1183), .Z(n476) );
  INV_X1 U153 ( .A(n1247), .ZN(n1226) );
  NAND2_X1 U156 ( .A1(n784), .A2(n1149), .ZN(n645) );
  INV_X1 U157 ( .A(n1475), .ZN(n1476) );
  NAND2_X1 U159 ( .A1(n1618), .A2(n1620), .ZN(n1687) );
  NAND2_X1 U160 ( .A1(n1750), .A2(n273), .ZN(n563) );
  NAND2_X1 U166 ( .A1(n41), .A2(n1159), .ZN(n196) );
  BUF_X2 U180 ( .A(n1351), .Z(n411) );
  NOR2_X2 U189 ( .A1(n562), .A2(n1271), .ZN(n1416) );
  NAND2_X1 U195 ( .A1(n1591), .A2(n1663), .ZN(n1589) );
  INV_X1 U204 ( .A(n1393), .ZN(n1311) );
  NOR2_X1 U213 ( .A1(n1429), .A2(n1428), .ZN(n1449) );
  BUF_X1 U220 ( .A(n1439), .Z(n250) );
  NOR2_X1 U225 ( .A1(n1461), .A2(n837), .ZN(n1739) );
  NAND2_X1 U227 ( .A1(n1435), .A2(n1434), .ZN(n1437) );
  BUF_X1 U233 ( .A(n269), .Z(n1575) );
  INV_X2 U245 ( .A(a[11]), .ZN(n978) );
  INV_X1 U250 ( .A(b[12]), .ZN(n120) );
  INV_X2 U255 ( .A(n1732), .ZN(n1247) );
  INV_X2 U264 ( .A(n994), .ZN(n1412) );
  INV_X1 U270 ( .A(n1521), .ZN(n163) );
  AND2_X2 U272 ( .A1(n903), .A2(a[15]), .ZN(n1668) );
  INV_X2 U273 ( .A(a[15]), .ZN(n1047) );
  INV_X2 U275 ( .A(a[19]), .ZN(n822) );
  NAND2_X2 U276 ( .A1(n1671), .A2(n1670), .ZN(\d[22] ) );
  AOI22_X2 U278 ( .A1(n431), .A2(n432), .B1(n422), .B2(n1661), .ZN(n1670) );
  NAND2_X2 U283 ( .A1(n198), .A2(n194), .ZN(n1671) );
  AOI22_X2 U286 ( .A1(n1265), .A2(n970), .B1(n971), .B2(n121), .ZN(n707) );
  NAND2_X2 U295 ( .A1(n231), .A2(n234), .ZN(n1287) );
  OAI21_X2 U311 ( .B1(n233), .B2(n850), .A(n1507), .ZN(n231) );
  NAND3_X2 U324 ( .A1(n262), .A2(n1404), .A3(n1402), .ZN(n1745) );
  NAND2_X2 U325 ( .A1(n1673), .A2(n1672), .ZN(n1119) );
  NAND3_X2 U334 ( .A1(n435), .A2(n729), .A3(n728), .ZN(n1672) );
  NAND2_X2 U335 ( .A1(n437), .A2(n1107), .ZN(n1673) );
  NAND3_X2 U337 ( .A1(n1336), .A2(n1495), .A3(n1334), .ZN(n188) );
  NAND2_X4 U339 ( .A1(n1298), .A2(n1299), .ZN(n1336) );
  NAND2_X2 U346 ( .A1(n369), .A2(n1156), .ZN(n464) );
  NAND2_X2 U347 ( .A1(n860), .A2(n863), .ZN(n1522) );
  NAND2_X2 U348 ( .A1(n1697), .A2(n861), .ZN(n860) );
  NAND2_X2 U351 ( .A1(n1007), .A2(n1006), .ZN(n1681) );
  NAND2_X2 U354 ( .A1(n938), .A2(n56), .ZN(n899) );
  XNOR2_X2 U357 ( .A(n541), .B(n51), .ZN(n921) );
  NAND2_X2 U361 ( .A1(n1572), .A2(n181), .ZN(n541) );
  INV_X2 U369 ( .A(n918), .ZN(n1298) );
  NAND3_X2 U377 ( .A1(n74), .A2(n1674), .A3(n1409), .ZN(\d[16]_BAR ) );
  AOI21_X2 U378 ( .B1(n1626), .B2(n1407), .A(n1406), .ZN(n1674) );
  OAI21_X2 U384 ( .B1(n1014), .B2(n545), .A(n1612), .ZN(n1017) );
  NAND2_X2 U385 ( .A1(n1461), .A2(n138), .ZN(n908) );
  AOI22_X2 U386 ( .A1(n1735), .A2(n913), .B1(n910), .B2(n909), .ZN(n1461) );
  AOI22_X2 U393 ( .A1(n1281), .A2(n765), .B1(n1420), .B2(n1280), .ZN(n1284) );
  NAND2_X2 U406 ( .A1(n211), .A2(n986), .ZN(n904) );
  NAND3_X2 U408 ( .A1(n905), .A2(n977), .A3(n976), .ZN(n211) );
  NAND3_X2 U409 ( .A1(n1484), .A2(n1675), .A3(n1482), .ZN(\d[15]_BAR ) );
  NOR2_X2 U410 ( .A1(n1479), .A2(n596), .ZN(n1675) );
  NAND2_X2 U411 ( .A1(n772), .A2(n773), .ZN(n213) );
  NAND2_X2 U416 ( .A1(n46), .A2(n866), .ZN(n772) );
  NAND3_X2 U419 ( .A1(n918), .A2(n920), .A3(n919), .ZN(n1337) );
  NAND2_X2 U420 ( .A1(n468), .A2(n989), .ZN(n769) );
  NOR2_X4 U424 ( .A1(n968), .A2(b[12]), .ZN(n468) );
  XNOR2_X2 U425 ( .A(n1511), .B(n1676), .ZN(n1012) );
  INV_X4 U427 ( .A(a[19]), .ZN(n1676) );
  NAND2_X2 U435 ( .A1(n843), .A2(n1089), .ZN(n875) );
  NOR2_X4 U439 ( .A1(n1194), .A2(n812), .ZN(n843) );
  NAND2_X2 U441 ( .A1(n1677), .A2(n1061), .ZN(n1090) );
  NAND2_X2 U442 ( .A1(n350), .A2(n1060), .ZN(n1677) );
  NAND2_X1 U444 ( .A1(n773), .A2(n772), .ZN(n1678) );
  INV_X4 U448 ( .A(n1093), .ZN(n873) );
  NOR2_X4 U455 ( .A1(n1093), .A2(n1094), .ZN(n754) );
  NAND2_X2 U459 ( .A1(n330), .A2(n110), .ZN(n1679) );
  NAND2_X2 U464 ( .A1(n330), .A2(n110), .ZN(n1030) );
  INV_X2 U467 ( .A(n866), .ZN(n865) );
  INV_X2 U469 ( .A(n1388), .ZN(n44) );
  NAND2_X2 U471 ( .A1(n986), .A2(n211), .ZN(n1680) );
  NAND2_X2 U478 ( .A1(n244), .A2(n243), .ZN(n270) );
  INV_X4 U484 ( .A(n406), .ZN(n158) );
  NOR2_X1 U486 ( .A1(a[10]), .A2(n798), .ZN(n1273) );
  NAND2_X1 U487 ( .A1(n893), .A2(n1657), .ZN(n1682) );
  INV_X2 U491 ( .A(n1310), .ZN(n1611) );
  INV_X2 U492 ( .A(n921), .ZN(n1715) );
  NOR2_X1 U493 ( .A1(n1387), .A2(n1386), .ZN(n322) );
  NAND2_X1 U495 ( .A1(n785), .A2(n1148), .ZN(n130) );
  INV_X4 U496 ( .A(n1051), .ZN(n687) );
  NAND2_X1 U497 ( .A1(n822), .A2(n820), .ZN(n821) );
  NAND2_X2 U505 ( .A1(n244), .A2(n243), .ZN(n1722) );
  INV_X4 U507 ( .A(n1701), .ZN(n1398) );
  AND2_X1 U508 ( .A1(n149), .A2(n150), .ZN(n1036) );
  INV_X1 U509 ( .A(n150), .ZN(n1618) );
  INV_X2 U512 ( .A(n263), .ZN(n539) );
  INV_X4 U514 ( .A(b[13]), .ZN(n1683) );
  INV_X4 U515 ( .A(b[13]), .ZN(n806) );
  NAND2_X4 U518 ( .A1(n718), .A2(n1473), .ZN(n135) );
  NAND2_X1 U521 ( .A1(n1604), .A2(n1603), .ZN(n1684) );
  NAND2_X2 U522 ( .A1(n1100), .A2(n1093), .ZN(n1101) );
  AND3_X1 U530 ( .A1(n1117), .A2(n1343), .A3(n1118), .ZN(n1685) );
  NAND2_X2 U534 ( .A1(n148), .A2(n1686), .ZN(\d[18] ) );
  NAND3_X1 U537 ( .A1(n809), .A2(n941), .A3(n959), .ZN(n1686) );
  OAI21_X2 U545 ( .B1(n1036), .B2(n685), .A(n1687), .ZN(n1464) );
  BUF_X4 U550 ( .A(n1625), .Z(n1688) );
  NAND2_X2 U552 ( .A1(n1351), .A2(n554), .ZN(n1355) );
  NAND2_X2 U554 ( .A1(n553), .A2(n1393), .ZN(n1351) );
  NOR2_X2 U556 ( .A1(n1216), .A2(n1689), .ZN(n528) );
  NOR3_X2 U563 ( .A1(n1215), .A2(n1221), .A3(n1214), .ZN(n1689) );
  NAND2_X4 U566 ( .A1(n371), .A2(n372), .ZN(n1349) );
  NAND3_X2 U575 ( .A1(n799), .A2(n1209), .A3(n965), .ZN(n738) );
  NAND3_X2 U579 ( .A1(n17), .A2(n133), .A3(n134), .ZN(n147) );
  NAND2_X2 U581 ( .A1(n189), .A2(n183), .ZN(n432) );
  NAND2_X2 U582 ( .A1(b[10]), .A2(n618), .ZN(n620) );
  NOR2_X2 U589 ( .A1(n551), .A2(n1220), .ZN(n600) );
  NAND2_X2 U590 ( .A1(n715), .A2(n714), .ZN(n551) );
  NAND2_X2 U596 ( .A1(n307), .A2(n1289), .ZN(n1744) );
  NAND2_X2 U599 ( .A1(n117), .A2(n1202), .ZN(n307) );
  NAND2_X2 U602 ( .A1(n1690), .A2(n128), .ZN(n513) );
  NAND2_X2 U607 ( .A1(n122), .A2(n1291), .ZN(n1690) );
  NOR2_X2 U621 ( .A1(n513), .A2(n1287), .ZN(n72) );
  NAND3_X2 U630 ( .A1(n1361), .A2(n204), .A3(n41), .ZN(n941) );
  NAND2_X2 U641 ( .A1(n1693), .A2(n1692), .ZN(n1577) );
  NAND2_X2 U649 ( .A1(n124), .A2(n163), .ZN(n1692) );
  NAND2_X2 U655 ( .A1(n1547), .A2(n1521), .ZN(n1693) );
  NAND2_X2 U662 ( .A1(n1613), .A2(n756), .ZN(n336) );
  NOR2_X4 U669 ( .A1(n989), .A2(n120), .ZN(n1613) );
  NAND2_X2 U672 ( .A1(n1121), .A2(n1120), .ZN(n1124) );
  NOR2_X2 U675 ( .A1(n1308), .A2(n1616), .ZN(n429) );
  XNOR2_X2 U676 ( .A(n1384), .B(n1382), .ZN(n1308) );
  INV_X2 U689 ( .A(n1373), .ZN(n1305) );
  NAND2_X2 U691 ( .A1(n1694), .A2(n1704), .ZN(n8) );
  NAND2_X2 U707 ( .A1(n1696), .A2(n1695), .ZN(n1694) );
  INV_X2 U712 ( .A(n404), .ZN(n1695) );
  INV_X2 U717 ( .A(n405), .ZN(n1696) );
  NAND2_X2 U718 ( .A1(n170), .A2(n172), .ZN(n1629) );
  NAND3_X2 U724 ( .A1(n171), .A2(n174), .A3(n245), .ZN(n170) );
  NAND2_X2 U725 ( .A1(n265), .A2(n62), .ZN(n174) );
  NAND2_X2 U726 ( .A1(n1726), .A2(n1585), .ZN(n265) );
  NAND2_X2 U728 ( .A1(n1361), .A2(n204), .ZN(n175) );
  NAND3_X2 U736 ( .A1(n1118), .A2(n1343), .A3(n1117), .ZN(n204) );
  NOR2_X4 U743 ( .A1(n1318), .A2(n37), .ZN(n1361) );
  NAND2_X1 U750 ( .A1(n1236), .A2(n1237), .ZN(n658) );
  AOI22_X2 U756 ( .A1(n1751), .A2(n859), .B1(n1522), .B2(n1226), .ZN(n1236) );
  NAND2_X1 U763 ( .A1(n65), .A2(n1412), .ZN(n1697) );
  OAI22_X2 U764 ( .A1(n1463), .A2(n1688), .B1(n1739), .B2(n1667), .ZN(\d[12] )
         );
  NAND2_X2 U766 ( .A1(n591), .A2(n822), .ZN(n1076) );
  NAND2_X2 U767 ( .A1(n1698), .A2(n956), .ZN(n1565) );
  NAND2_X2 U788 ( .A1(n1312), .A2(n35), .ZN(n1698) );
  NAND2_X2 U789 ( .A1(n1153), .A2(n751), .ZN(n1559) );
  NAND2_X2 U792 ( .A1(n1700), .A2(n1699), .ZN(n278) );
  INV_X2 U793 ( .A(n742), .ZN(n1699) );
  AOI21_X2 U794 ( .B1(n1079), .B2(n1080), .A(n1078), .ZN(n742) );
  NAND2_X2 U795 ( .A1(n569), .A2(n567), .ZN(n1700) );
  NAND2_X2 U796 ( .A1(n1719), .A2(n1617), .ZN(n1701) );
  NOR2_X2 U804 ( .A1(n1355), .A2(n1309), .ZN(n1719) );
  NOR2_X4 U809 ( .A1(n1703), .A2(n1702), .ZN(n1039) );
  INV_X2 U812 ( .A(n822), .ZN(n1702) );
  INV_X4 U815 ( .A(n394), .ZN(n1703) );
  AOI21_X2 U822 ( .B1(n1130), .B2(a[12]), .A(n808), .ZN(n624) );
  NAND2_X1 U829 ( .A1(n591), .A2(n991), .ZN(n579) );
  NAND3_X1 U836 ( .A1(n552), .A2(n1487), .A3(n1466), .ZN(n1471) );
  NAND2_X2 U843 ( .A1(n1076), .A2(n1077), .ZN(n1078) );
  INV_X4 U853 ( .A(n281), .ZN(n352) );
  NAND3_X2 U864 ( .A1(n351), .A2(n354), .A3(n353), .ZN(n281) );
  NAND2_X2 U871 ( .A1(n722), .A2(n520), .ZN(n1539) );
  NAND2_X2 U872 ( .A1(n1580), .A2(n1579), .ZN(n722) );
  NAND2_X2 U873 ( .A1(n405), .A2(n404), .ZN(n1704) );
  NOR2_X2 U875 ( .A1(n1705), .A2(n844), .ZN(n261) );
  NOR3_X2 U881 ( .A1(n255), .A2(n514), .A3(n254), .ZN(n1705) );
  NAND2_X4 U882 ( .A1(n888), .A2(n1459), .ZN(n359) );
  NAND2_X2 U883 ( .A1(n1679), .A2(n838), .ZN(n1459) );
  NAND2_X4 U884 ( .A1(n1172), .A2(n1706), .ZN(n364) );
  NAND2_X2 U886 ( .A1(n1170), .A2(n589), .ZN(n1706) );
  NOR2_X2 U890 ( .A1(n804), .A2(n897), .ZN(n1487) );
  NAND2_X2 U891 ( .A1(n169), .A2(n167), .ZN(n1439) );
  NAND2_X2 U901 ( .A1(n1284), .A2(n1418), .ZN(n1752) );
  NOR2_X4 U902 ( .A1(n1707), .A2(n1135), .ZN(n655) );
  NAND2_X2 U904 ( .A1(n1127), .A2(n1126), .ZN(n1707) );
  NAND2_X2 U905 ( .A1(n722), .A2(n520), .ZN(n68) );
  NOR2_X2 U908 ( .A1(n104), .A2(n1125), .ZN(n706) );
  NAND2_X2 U916 ( .A1(n1708), .A2(n1525), .ZN(n1004) );
  NAND2_X2 U917 ( .A1(n689), .A2(n1047), .ZN(n1708) );
  NAND2_X1 U920 ( .A1(n673), .A2(n674), .ZN(n1163) );
  NAND2_X1 U924 ( .A1(n527), .A2(n219), .ZN(n218) );
  NAND2_X1 U931 ( .A1(n1136), .A2(n625), .ZN(n221) );
  INV_X2 U935 ( .A(n467), .ZN(n1152) );
  AOI22_X2 U936 ( .A1(n680), .A2(n857), .B1(n855), .B2(n1067), .ZN(n1709) );
  NAND2_X1 U937 ( .A1(n1495), .A2(n1334), .ZN(n1335) );
  INV_X1 U945 ( .A(n1495), .ZN(n1322) );
  AOI22_X1 U953 ( .A1(n1477), .A2(n262), .B1(n1476), .B2(n851), .ZN(n1478) );
  AOI21_X2 U959 ( .B1(n752), .B2(n735), .A(n1081), .ZN(n1710) );
  NOR2_X4 U969 ( .A1(n1050), .A2(n752), .ZN(n1081) );
  INV_X2 U990 ( .A(n115), .ZN(n1635) );
  NAND2_X1 U995 ( .A1(n907), .A2(n1623), .ZN(n1713) );
  NAND2_X2 U996 ( .A1(n1713), .A2(n1714), .ZN(n176) );
  INV_X2 U1014 ( .A(n335), .ZN(n1595) );
  INV_X1 U1017 ( .A(n1231), .ZN(n241) );
  NAND2_X1 U1020 ( .A1(n928), .A2(n489), .ZN(n983) );
  XNOR2_X1 U1021 ( .A(n489), .B(n636), .ZN(n565) );
  INV_X2 U1022 ( .A(n1727), .ZN(n545) );
  NAND2_X2 U1027 ( .A1(n871), .A2(n870), .ZN(n62) );
  NAND2_X1 U1033 ( .A1(n921), .A2(n1305), .ZN(n1717) );
  NAND2_X2 U1039 ( .A1(n1715), .A2(n1716), .ZN(n1718) );
  NAND2_X2 U1041 ( .A1(n1717), .A2(n1718), .ZN(n918) );
  INV_X1 U1048 ( .A(n1305), .ZN(n1716) );
  INV_X2 U1060 ( .A(n1752), .ZN(n379) );
  NAND3_X2 U1079 ( .A1(n1293), .A2(n89), .A3(n628), .ZN(n1720) );
  NAND3_X1 U1082 ( .A1(n1293), .A2(n89), .A3(n628), .ZN(n1633) );
  XNOR2_X1 U1083 ( .A(n790), .B(n671), .ZN(n789) );
  NAND2_X1 U1088 ( .A1(n751), .A2(n755), .ZN(n641) );
  NAND2_X1 U1093 ( .A1(n412), .A2(n994), .ZN(n861) );
  NAND2_X2 U1095 ( .A1(n1719), .A2(n1617), .ZN(n1721) );
  INV_X1 U1097 ( .A(n8), .ZN(n543) );
  NAND2_X1 U1103 ( .A1(n808), .A2(n1723), .ZN(n1724) );
  NAND2_X2 U1112 ( .A1(n472), .A2(n1412), .ZN(n1725) );
  NAND2_X2 U1113 ( .A1(n1724), .A2(n1725), .ZN(n1254) );
  INV_X1 U1120 ( .A(n1412), .ZN(n1723) );
  NOR2_X4 U1128 ( .A1(n845), .A2(n822), .ZN(n1038) );
  AOI21_X1 U1130 ( .B1(n1332), .B2(n175), .A(n1329), .ZN(n1330) );
  AOI21_X1 U1137 ( .B1(n1046), .B2(b[8]), .A(n1045), .ZN(n735) );
  NAND2_X2 U1143 ( .A1(n268), .A2(n1108), .ZN(n1726) );
  NAND2_X2 U1145 ( .A1(n1217), .A2(n1231), .ZN(n1230) );
  NOR2_X2 U1153 ( .A1(n528), .A2(n1232), .ZN(n1231) );
  NAND2_X2 U1154 ( .A1(n1212), .A2(n1213), .ZN(n1727) );
  NAND2_X2 U1155 ( .A1(n1728), .A2(n1515), .ZN(n1258) );
  NAND2_X2 U1158 ( .A1(n1513), .A2(a[11]), .ZN(n1728) );
  INV_X4 U1169 ( .A(n1729), .ZN(n96) );
  NOR2_X2 U1178 ( .A1(n601), .A2(n1632), .ZN(n1729) );
  NAND3_X2 U1185 ( .A1(n807), .A2(n994), .A3(b[14]), .ZN(n1601) );
  NAND2_X2 U1187 ( .A1(n1296), .A2(n8), .ZN(n775) );
  AOI22_X2 U1188 ( .A1(n1749), .A2(n1187), .B1(n1186), .B2(n406), .ZN(n1296)
         );
  NAND2_X2 U1196 ( .A1(n937), .A2(a[13]), .ZN(n1011) );
  NAND2_X4 U1197 ( .A1(n1511), .A2(n962), .ZN(n104) );
  NOR2_X2 U1205 ( .A1(n968), .A2(n965), .ZN(n962) );
  BUF_X4 U1217 ( .A(n1403), .Z(n1730) );
  NAND2_X2 U1226 ( .A1(n1430), .A2(n1425), .ZN(n484) );
  AND2_X2 U1228 ( .A1(n1617), .A2(n1310), .ZN(n1735) );
  INV_X2 U1237 ( .A(a[8]), .ZN(n1733) );
  AOI21_X2 U1244 ( .B1(n937), .B2(n18), .A(n1733), .ZN(n1732) );
  INV_X4 U1258 ( .A(n1734), .ZN(n1756) );
  NAND2_X2 U1267 ( .A1(n863), .A2(n860), .ZN(n1734) );
  NAND2_X2 U1269 ( .A1(n234), .A2(n231), .ZN(n1521) );
  INV_X2 U1272 ( .A(n1275), .ZN(n1278) );
  NAND2_X2 U1274 ( .A1(n1737), .A2(n1736), .ZN(n1275) );
  NAND2_X2 U1288 ( .A1(n845), .A2(n1412), .ZN(n1736) );
  NAND2_X2 U1290 ( .A1(n1270), .A2(n994), .ZN(n1737) );
  NAND3_X1 U1292 ( .A1(n863), .A2(n860), .A3(n1247), .ZN(n859) );
  NAND2_X2 U1313 ( .A1(n1225), .A2(n757), .ZN(n863) );
  NOR2_X4 U1314 ( .A1(n984), .A2(n1738), .ZN(n1021) );
  NAND3_X2 U1318 ( .A1(n1741), .A2(n982), .A3(n1740), .ZN(n1738) );
  NAND2_X2 U1325 ( .A1(n1569), .A2(a[12]), .ZN(n1740) );
  NAND2_X2 U1327 ( .A1(n988), .A2(n820), .ZN(n1741) );
  NAND2_X2 U1328 ( .A1(n68), .A2(n67), .ZN(n71) );
  NAND2_X2 U1332 ( .A1(n1628), .A2(n1088), .ZN(n67) );
  NAND2_X2 U1344 ( .A1(n1207), .A2(n1208), .ZN(n1222) );
  NAND2_X2 U1349 ( .A1(n1205), .A2(n1206), .ZN(n1207) );
  NAND2_X2 U1366 ( .A1(n723), .A2(n539), .ZN(n1640) );
  INV_X2 U1367 ( .A(n1742), .ZN(n1641) );
  NAND2_X2 U1371 ( .A1(n916), .A2(n271), .ZN(n1742) );
  INV_X4 U1377 ( .A(b[14]), .ZN(n1022) );
  NAND2_X2 U1378 ( .A1(n1744), .A2(n1743), .ZN(n122) );
  INV_X2 U1386 ( .A(n1288), .ZN(n1743) );
  NAND3_X2 U1387 ( .A1(n923), .A2(n1745), .A3(n1405), .ZN(n1406) );
  BUF_X4 U1398 ( .A(n1509), .Z(n1746) );
  INV_X2 U1404 ( .A(n301), .ZN(n677) );
  NAND2_X2 U1418 ( .A1(n1505), .A2(n1747), .ZN(n301) );
  NAND2_X1 U1426 ( .A1(n203), .A2(n1072), .ZN(n1747) );
  INV_X4 U1448 ( .A(n1179), .ZN(n1748) );
  NOR3_X2 U1455 ( .A1(n1096), .A2(n1097), .A3(n1095), .ZN(n1099) );
  NAND2_X2 U1456 ( .A1(n158), .A2(n157), .ZN(n1749) );
  NAND2_X2 U1472 ( .A1(n1344), .A2(n1503), .ZN(n1339) );
  NOR3_X2 U1484 ( .A1(n1335), .A2(n2), .A3(n638), .ZN(n1344) );
  NAND2_X2 U1490 ( .A1(n1517), .A2(n943), .ZN(n942) );
  XNOR2_X2 U1499 ( .A(n808), .B(n1750), .ZN(n1225) );
  INV_X2 U1504 ( .A(a[10]), .ZN(n1750) );
  NAND2_X2 U1505 ( .A1(n853), .A2(n864), .ZN(n1751) );
  NAND2_X2 U1506 ( .A1(n317), .A2(n1752), .ZN(n1293) );
  NOR2_X2 U1513 ( .A1(n1355), .A2(n1309), .ZN(n317) );
  NAND3_X2 U1517 ( .A1(n70), .A2(n1539), .A3(n67), .ZN(n721) );
  NAND2_X2 U1518 ( .A1(n374), .A2(n373), .ZN(n70) );
  NAND2_X2 U1527 ( .A1(n1756), .A2(n1226), .ZN(n80) );
  AOI22_X2 U1529 ( .A1(n561), .A2(n746), .B1(n1753), .B2(n1200), .ZN(n124) );
  NAND2_X2 U1534 ( .A1(n161), .A2(n13), .ZN(n1753) );
  NAND2_X2 U1536 ( .A1(n90), .A2(n531), .ZN(n88) );
  NAND2_X2 U1546 ( .A1(n950), .A2(n281), .ZN(n90) );
  NAND2_X2 U1556 ( .A1(n1400), .A2(n613), .ZN(n1364) );
  NAND2_X2 U1558 ( .A1(n1554), .A2(n306), .ZN(n1400) );
  NAND2_X2 U1559 ( .A1(n82), .A2(n1754), .ZN(n1276) );
  NAND2_X2 U1560 ( .A1(n257), .A2(a[8]), .ZN(n1754) );
  NOR2_X2 U1561 ( .A1(n472), .A2(n1130), .ZN(n471) );
  NOR2_X2 U1562 ( .A1(n1755), .A2(n1401), .ZN(n596) );
  INV_X2 U1563 ( .A(n1481), .ZN(n1755) );
  NOR2_X2 U1564 ( .A1(n262), .A2(n1475), .ZN(n1481) );
  INV_X4 U1565 ( .A(n168), .ZN(n461) );
  INV_X4 U1566 ( .A(n1349), .ZN(n1540) );
  INV_X2 U1161 ( .A(a[25]), .ZN(n952) );
  OAI21_X1 U101 ( .B1(n1444), .B2(n1446), .A(n1757), .ZN(\d[3] ) );
  AOI22_X1 U102 ( .A1(n1448), .A2(n1449), .B1(n1444), .B2(n1758), .ZN(n1757)
         );
  INV_X1 U135 ( .A(n1445), .ZN(n1758) );
  OAI211_X1 U140 ( .C1(n138), .C2(n837), .A(n613), .B(n1759), .ZN(n1667) );
  OR2_X1 U209 ( .A1(n898), .A2(n897), .ZN(n1759) );
  INV_X1 U228 ( .A(n1393), .ZN(n1760) );
  NOR2_X2 U229 ( .A1(n1760), .A2(n610), .ZN(n23) );
  INV_X1 U240 ( .A(n1761), .ZN(n1564) );
  AOI22_X1 U243 ( .A1(n1540), .A2(n1503), .B1(n1349), .B2(n1348), .ZN(n1761)
         );
  AND2_X2 U246 ( .A1(n16), .A2(n17), .ZN(n1319) );
  INV_X1 U247 ( .A(n1113), .ZN(n1762) );
  NAND2_X2 U274 ( .A1(n1762), .A2(n1109), .ZN(n598) );
  INV_X1 U400 ( .A(n1763), .ZN(n1714) );
  NOR2_X2 U404 ( .A1(n907), .A2(n1623), .ZN(n1763) );
  OAI21_X1 U494 ( .B1(a[11]), .B2(n776), .A(n1764), .ZN(n1274) );
  NAND2_X1 U498 ( .A1(n947), .A2(a[11]), .ZN(n1764) );
  OAI21_X1 U633 ( .B1(n1376), .B2(n55), .A(n1765), .ZN(n1306) );
  NAND2_X1 U637 ( .A1(n55), .A2(n732), .ZN(n1765) );
  INV_X1 U640 ( .A(a[8]), .ZN(n283) );
  AND2_X1 U715 ( .A1(a[8]), .A2(b[10]), .ZN(n636) );
  OR2_X2 U790 ( .A1(n591), .A2(a[11]), .ZN(n339) );
  OR2_X2 U791 ( .A1(n969), .A2(n887), .ZN(n1658) );
  AND2_X2 U892 ( .A1(n38), .A2(a[25]), .ZN(n603) );
endmodule

