library verilog;
use verilog.vl_types.all;
entity CLKBUF_X1_func is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end CLKBUF_X1_func;
