library verilog;
use verilog.vl_types.all;
entity MUX2_X1_func is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        S               : in     vl_logic;
        Z               : out    vl_logic
    );
end MUX2_X1_func;
