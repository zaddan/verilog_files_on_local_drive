//*** remember that I have removed the dummy and commented out everything about it
module conf_int_mul__noFF__arch_agnos_OP_BITWIDTH18_DATA_PATH_BITWIDTH26__acc ( clk, 
        racc, rapx, a, b, \d[40] , \d[39] , \d[36] , \d[34] , \d[32] , \d[29] , 
        \d[25] , \d[23] , \d[11] , \d[7] , \d[6] , \d[5] , \d[4] , \d[3] , 
        \d[2] , \d[1] , \d[0] , \d[37]_BAR , \d[30]_BAR , \d[24]_BAR , 
        \d[21]_BAR , \d[20]_BAR , \d[14]_BAR , \d[9]_BAR , \d[8]_BAR , \d[28] , 
        \d[27]_BAR , \d[31]_BAR , \d[17] , \d[13]_BAR , \d[35]_BAR , \d[19] , 
        \d[22]_BAR , \d[15]_BAR , \d[18] , \d[10]_BAR , \d[16]_BAR , \d[33] , 
        \d[38]_BAR , \d[12]_BAR , \d[26]  );
  input [25:0] a;
  input [14:0] b;
  input clk, racc, rapx;
  output \d[40] , \d[39] , \d[36] , \d[34] , \d[32] , \d[29] , \d[25] ,
         \d[23] , \d[11] , \d[7] , \d[6] , \d[5] , \d[4] , \d[3] , \d[2] ,
         \d[1] , \d[0] , \d[37]_BAR , \d[30]_BAR , \d[24]_BAR , \d[21]_BAR ,
         \d[20]_BAR , \d[14]_BAR , \d[9]_BAR , \d[8]_BAR , \d[28] ,
         \d[27]_BAR , \d[31]_BAR , \d[17] , \d[13]_BAR , \d[35]_BAR , \d[19] ,
         \d[22]_BAR , \d[15]_BAR , \d[18] , \d[10]_BAR , \d[16]_BAR , \d[33] ,
         \d[38]_BAR , \d[12]_BAR , \d[26] ;
  wire   n1, n2, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n107, n109,
         n110, n111, n115, n116, n117, n118, n119, n121, n123, n124, n127,
         n128, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n150, n151,
         n152, n155, n156, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n184, n185, n186, n187, n188, n189,
         n191, n192, n193, n194, n196, n197, n198, n199, n200, n201, n203,
         n204, n205, n206, n207, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n224, n225, n226, n227, n228,
         n230, n231, n232, n233, n234, n235, n236, n237, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n322,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n360, n362, n363, n364, n365, n366, n367, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n409, n410, n411, n412, n413, n414, n415, n418, n419,
         n420, n421, n422, n424, n425, n426, n427, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n469, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n670, n671, n672, n673, n674, n675, n677, n678, n679,
         n680, n681, n682, n683, n684, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n740, n741, n742, n743, n744, n746, n748, n749, n750, n751,
         n752, n753, n756, n757, n758, n759, n760, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n861,
         n862, n863, n864, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n911, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n954, n955, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1012, n1013, n1014, n1015,
         n1016, n1019, n1021, n1022, n1023, n1024, n1025, n1029, n1030, n1033,
         n1034, n1036, n1037, n1038, n1039, n1040, n1041, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1113, n1116, n1117, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1179, n1180, n1181,
         n1182, n1184, n1185, n1186, n1187, n1188, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1204, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1219, n1220,
         n1221, n1222, n1223, n1224, n1226, n1227, n1228, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1250, n1251, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1342, n1343, n1344, n1346, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1392, n1393, n1395, n1396, n1397, n1398, n1399, n1400, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1512, n1513, n1514, n1517, n1518, n1519, n1520, n1521, n1524,
         n1525, n1528, n1529, n1530, n1531, n1532, n1533, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1589, n1590, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1699, n1701, n1702, n1703, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1715, n1716, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1756, n1757, n1758,
         n1759, n1760, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1779, n1780,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1795, n1796,
         n1799, n1801, n1802, n1803, n1804, n1805, n1808, n1809, n1810, n1811,
         n1812, n1814, n1815, n1816, n1817, n1818, n1819, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1924, n1925, n1926, n1927, n1928, n1930, n1931, n1932,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1942, n1943, n1944,
         n1947, n1948, n1949, n1952, n1953, n1954, n1955, n1956, n1957, n1959,
         n1960, n1961, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2022, n2023, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2053, n2054,
         n2055, n2057, n2058, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2120, n2122,
         n2123, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2151, n2152, n2153, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2269, n2270, n2271, n2272, n2273, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2373, n2374, n2375, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2392, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2404, n2405, n2407, n2408, n2410, n2411, n2412, n2413,
         n2414, n2415, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2611, n2612, n2613, n2614,
         n2615, n2616, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2760, n2761, n2762, n2764, n2765, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2796, n2797, n2798, n2800,
         n2801, n2802, n2803, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2880, n2881, n2882, n2883, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2933, n2934, n2935, n2936, n2937, n2938,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3208, n3209, n3210, n3211, n3212, n3215, n3216, n3217,
         n3220, n3221, n3222, n3223, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3441, n3442, n3443, n3444, n3446, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3471, n3472, n3473,
         n3474, n3475, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3500, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3774, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4146, n4147, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4161, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4244, n4245;

  BUF_X4 U1 ( .A(n3494), .Z(n25) );
  BUF_X4 U2 ( .A(n3763), .Z(n43) );
  INV_X4 U4 ( .A(n1603), .ZN(n3990) );
  INV_X4 U6 ( .A(n31), .ZN(n771) );
  NOR2_X2 U8 ( .A1(n2448), .A2(n2447), .ZN(n1870) );
  BUF_X4 U11 ( .A(n3023), .Z(n34) );
  INV_X2 U16 ( .A(a[3]), .ZN(n3534) );
  INV_X1 U18 ( .A(n1318), .ZN(n3897) );
  NAND2_X2 U23 ( .A1(n2812), .A2(n872), .ZN(n1163) );
  NAND2_X4 U24 ( .A1(n962), .A2(n961), .ZN(n2812) );
  NAND2_X2 U27 ( .A1(n1537), .A2(n2816), .ZN(n227) );
  INV_X8 U28 ( .A(n3475), .ZN(n58) );
  NAND2_X2 U29 ( .A1(n4023), .A2(n1508), .ZN(n3946) );
  NAND2_X2 U30 ( .A1(n3735), .A2(n3734), .ZN(n4023) );
  OAI21_X2 U32 ( .B1(n2), .B2(n1), .A(n1699), .ZN(n243) );
  NAND2_X2 U33 ( .A1(n1555), .A2(n57), .ZN(n1) );
  NAND3_X2 U36 ( .A1(n1940), .A2(n1710), .A3(n4169), .ZN(n305) );
  OAI21_X2 U37 ( .B1(n1830), .B2(n3022), .A(n3021), .ZN(n1940) );
  NAND3_X2 U40 ( .A1(n2341), .A2(n3895), .A3(n3891), .ZN(n3969) );
  INV_X4 U43 ( .A(n934), .ZN(n139) );
  NAND2_X2 U44 ( .A1(n4), .A2(n545), .ZN(n544) );
  NAND2_X2 U45 ( .A1(n4093), .A2(n78), .ZN(n4) );
  NOR2_X2 U46 ( .A1(n3667), .A2(n855), .ZN(n3656) );
  NOR2_X2 U47 ( .A1(n854), .A2(n3852), .ZN(n3667) );
  NAND2_X2 U49 ( .A1(n541), .A2(n543), .ZN(n324) );
  NAND3_X2 U58 ( .A1(n2281), .A2(n1701), .A3(n1232), .ZN(n3021) );
  NAND2_X2 U59 ( .A1(n7), .A2(n8), .ZN(n116) );
  NAND2_X2 U60 ( .A1(n144), .A2(n2922), .ZN(n7) );
  NAND3_X2 U61 ( .A1(n145), .A2(n1877), .A3(n1876), .ZN(n8) );
  NAND2_X2 U62 ( .A1(n194), .A2(n2358), .ZN(n2294) );
  INV_X2 U65 ( .A(n243), .ZN(n9) );
  BUF_X4 U67 ( .A(n3174), .Z(n10) );
  NAND2_X2 U68 ( .A1(n12), .A2(n11), .ZN(n2943) );
  NAND2_X2 U70 ( .A1(n1466), .A2(n1465), .ZN(n12) );
  NAND2_X2 U73 ( .A1(n13), .A2(n1475), .ZN(n102) );
  NAND2_X2 U74 ( .A1(n1582), .A2(n1581), .ZN(n13) );
  NAND2_X2 U75 ( .A1(n898), .A2(n2977), .ZN(n897) );
  AOI21_X1 U77 ( .B1(n3475), .B2(n249), .A(n3010), .ZN(n959) );
  NAND2_X2 U78 ( .A1(n1281), .A2(n2282), .ZN(n3020) );
  NAND2_X2 U79 ( .A1(n1232), .A2(n1701), .ZN(n1281) );
  INV_X1 U82 ( .A(a[14]), .ZN(n2239) );
  NOR2_X1 U83 ( .A1(n2938), .A2(n982), .ZN(n981) );
  NAND2_X1 U84 ( .A1(n84), .A2(n3407), .ZN(n636) );
  INV_X1 U85 ( .A(a[13]), .ZN(n2077) );
  NAND2_X1 U86 ( .A1(n86), .A2(n2057), .ZN(n2260) );
  INV_X1 U87 ( .A(n3162), .ZN(n1009) );
  NAND2_X1 U88 ( .A1(n1995), .A2(n1996), .ZN(n1722) );
  NAND2_X1 U89 ( .A1(n1862), .A2(n2258), .ZN(n493) );
  NAND2_X1 U90 ( .A1(n2044), .A2(n1658), .ZN(n1857) );
  INV_X4 U92 ( .A(n2506), .ZN(n3498) );
  NOR2_X1 U95 ( .A1(n942), .A2(n1870), .ZN(n939) );
  NAND2_X1 U96 ( .A1(n1068), .A2(n1067), .ZN(n1066) );
  NAND3_X1 U97 ( .A1(n1873), .A2(n2252), .A3(n2504), .ZN(n1871) );
  NAND2_X1 U98 ( .A1(n703), .A2(n702), .ZN(n3033) );
  INV_X1 U101 ( .A(n3316), .ZN(n3317) );
  NAND3_X1 U102 ( .A1(n2364), .A2(n1096), .A3(n2363), .ZN(n1094) );
  NAND2_X1 U104 ( .A1(n2601), .A2(n2600), .ZN(n731) );
  INV_X1 U105 ( .A(n789), .ZN(n788) );
  NAND2_X1 U106 ( .A1(n3413), .A2(n3431), .ZN(n422) );
  NOR2_X1 U107 ( .A1(n3432), .A2(n452), .ZN(n518) );
  NAND2_X1 U108 ( .A1(n66), .A2(n3559), .ZN(n3369) );
  NOR2_X1 U110 ( .A1(n1745), .A2(n3947), .ZN(n1619) );
  NAND3_X1 U112 ( .A1(n3854), .A2(n3620), .A3(n3722), .ZN(n3637) );
  OR2_X4 U113 ( .A1(n3576), .A2(n3575), .ZN(n14) );
  INV_X1 U114 ( .A(n3172), .ZN(n2317) );
  AND2_X4 U118 ( .A1(n1815), .A2(n1814), .ZN(n18) );
  OR2_X4 U119 ( .A1(n267), .A2(n1752), .ZN(n19) );
  AND2_X2 U120 ( .A1(n1978), .A2(n1977), .ZN(n20) );
  AND2_X4 U121 ( .A1(n3190), .A2(n3184), .ZN(n21) );
  AND2_X4 U124 ( .A1(n674), .A2(n1395), .ZN(n22) );
  NOR2_X1 U127 ( .A1(n2155), .A2(n1236), .ZN(n1070) );
  INV_X1 U128 ( .A(n35), .ZN(n2475) );
  INV_X1 U129 ( .A(n3377), .ZN(n3378) );
  AND2_X4 U130 ( .A1(n3075), .A2(n3076), .ZN(n24) );
  INV_X4 U131 ( .A(n3139), .ZN(n56) );
  INV_X1 U132 ( .A(n3380), .ZN(n1878) );
  INV_X1 U133 ( .A(a[11]), .ZN(n3118) );
  INV_X1 U135 ( .A(n3906), .ZN(n3833) );
  NOR2_X1 U136 ( .A1(n3984), .A2(n4207), .ZN(n3903) );
  NAND2_X1 U141 ( .A1(n3737), .A2(n4032), .ZN(n3569) );
  NAND2_X1 U142 ( .A1(n1464), .A2(n1844), .ZN(n1321) );
  OR2_X2 U143 ( .A1(n87), .A2(a[24]), .ZN(n174) );
  NAND3_X1 U144 ( .A1(n1025), .A2(n461), .A3(n3330), .ZN(n3331) );
  NAND2_X2 U145 ( .A1(n427), .A2(n1337), .ZN(n426) );
  NAND3_X1 U146 ( .A1(n38), .A2(n4048), .A3(n36), .ZN(n35) );
  NOR2_X1 U148 ( .A1(n30), .A2(n29), .ZN(n2312) );
  NOR2_X1 U149 ( .A1(n3080), .A2(a[17]), .ZN(n29) );
  NOR2_X1 U150 ( .A1(n1303), .A2(n3124), .ZN(n30) );
  NAND3_X1 U151 ( .A1(n3563), .A2(n3926), .A3(n3562), .ZN(n3932) );
  NAND4_X1 U152 ( .A1(n600), .A2(n1172), .A3(n1171), .A4(n1170), .ZN(n1536) );
  NAND4_X1 U153 ( .A1(n318), .A2(n2161), .A3(n426), .A4(n317), .ZN(n314) );
  INV_X2 U156 ( .A(n2146), .ZN(n31) );
  NAND2_X1 U158 ( .A1(n1337), .A2(n3069), .ZN(n32) );
  NAND2_X1 U160 ( .A1(n1928), .A2(n45), .ZN(n279) );
  AOI22_X1 U161 ( .A1(n3034), .A2(n56), .B1(n249), .B2(a[8]), .ZN(n278) );
  NAND2_X1 U162 ( .A1(n2737), .A2(n37), .ZN(n36) );
  INV_X1 U163 ( .A(n3124), .ZN(n37) );
  NAND2_X1 U164 ( .A1(n2736), .A2(n3124), .ZN(n38) );
  AND2_X2 U166 ( .A1(n3058), .A2(n3057), .ZN(n1197) );
  NAND2_X1 U168 ( .A1(n46), .A2(n45), .ZN(n44) );
  INV_X1 U170 ( .A(n3329), .ZN(n46) );
  NAND2_X1 U171 ( .A1(n2315), .A2(a[23]), .ZN(n47) );
  NAND2_X1 U173 ( .A1(n918), .A2(n2836), .ZN(n2837) );
  NAND3_X1 U174 ( .A1(n48), .A2(n889), .A3(n888), .ZN(n3900) );
  INV_X2 U175 ( .A(n891), .ZN(n48) );
  NAND2_X1 U176 ( .A1(n3893), .A2(n3895), .ZN(n891) );
  NOR3_X2 U177 ( .A1(n450), .A2(n4052), .A3(n2558), .ZN(n3241) );
  NAND2_X2 U178 ( .A1(n1872), .A2(n1871), .ZN(n1541) );
  INV_X1 U180 ( .A(n3164), .ZN(n2235) );
  INV_X1 U181 ( .A(n714), .ZN(n3386) );
  OR2_X4 U182 ( .A1(n3285), .A2(n3284), .ZN(n51) );
  INV_X1 U185 ( .A(n3947), .ZN(n3738) );
  NAND2_X4 U186 ( .A1(n274), .A2(n273), .ZN(n2966) );
  INV_X2 U188 ( .A(n4004), .ZN(n3954) );
  INV_X2 U189 ( .A(n2603), .ZN(n2604) );
  INV_X1 U190 ( .A(n1371), .ZN(n854) );
  NOR2_X4 U192 ( .A1(n3145), .A2(n3138), .ZN(n3154) );
  NAND2_X1 U193 ( .A1(n4003), .A2(n3978), .ZN(n1305) );
  NOR3_X1 U194 ( .A1(n4031), .A2(n3856), .A3(n3665), .ZN(n3671) );
  INV_X2 U195 ( .A(n3913), .ZN(n647) );
  INV_X2 U196 ( .A(n4005), .ZN(n1508) );
  AND2_X1 U198 ( .A1(n3988), .A2(n3987), .ZN(n472) );
  OR2_X1 U199 ( .A1(n3912), .A2(n1787), .ZN(n457) );
  INV_X2 U201 ( .A(n3617), .ZN(n3854) );
  NOR2_X2 U202 ( .A1(n2774), .A2(n2775), .ZN(n3374) );
  OR2_X1 U204 ( .A1(n2667), .A2(n2668), .ZN(n2669) );
  OAI21_X1 U206 ( .B1(n3401), .B2(n3402), .A(n3403), .ZN(n642) );
  AND2_X1 U207 ( .A1(n878), .A2(n874), .ZN(n473) );
  INV_X2 U208 ( .A(n2631), .ZN(n79) );
  NAND2_X2 U210 ( .A1(n2201), .A2(n2079), .ZN(n2265) );
  NOR2_X2 U212 ( .A1(n1819), .A2(n1822), .ZN(n2546) );
  INV_X4 U215 ( .A(n2620), .ZN(n53) );
  INV_X4 U217 ( .A(n1377), .ZN(n84) );
  NAND2_X2 U218 ( .A1(n3427), .A2(a[11]), .ZN(n2221) );
  INV_X2 U219 ( .A(n2989), .ZN(n89) );
  OR2_X2 U220 ( .A1(n3208), .A2(n2079), .ZN(n476) );
  AND2_X1 U221 ( .A1(n1835), .A2(a[7]), .ZN(n448) );
  INV_X4 U222 ( .A(n2924), .ZN(n92) );
  INV_X2 U223 ( .A(n1221), .ZN(n90) );
  INV_X2 U224 ( .A(n3202), .ZN(n94) );
  INV_X4 U225 ( .A(n2228), .ZN(n93) );
  INV_X4 U226 ( .A(n97), .ZN(n54) );
  INV_X2 U227 ( .A(a[18]), .ZN(n2442) );
  INV_X4 U228 ( .A(n3128), .ZN(n55) );
  INV_X4 U229 ( .A(a[14]), .ZN(n2438) );
  INV_X4 U230 ( .A(n3176), .ZN(n57) );
  AOI22_X1 U232 ( .A1(n3671), .A2(n3670), .B1(n3669), .B2(n3668), .ZN(n3672)
         );
  OAI21_X1 U233 ( .B1(n3827), .B2(n3904), .A(n3828), .ZN(n3795) );
  NAND2_X1 U235 ( .A1(n3878), .A2(n3877), .ZN(n3879) );
  INV_X1 U238 ( .A(n3949), .ZN(n3950) );
  INV_X2 U239 ( .A(n3928), .ZN(n3923) );
  NOR2_X1 U240 ( .A1(n3965), .A2(n3964), .ZN(n3976) );
  NAND2_X2 U241 ( .A1(n1620), .A2(n1619), .ZN(n4011) );
  INV_X2 U242 ( .A(n3635), .ZN(n3636) );
  AND2_X1 U243 ( .A1(n3912), .A2(n216), .ZN(n3914) );
  OR2_X2 U244 ( .A1(n3906), .A2(n3904), .ZN(n298) );
  NAND2_X2 U247 ( .A1(n3620), .A2(n3722), .ZN(n1846) );
  BUF_X4 U248 ( .A(n3911), .Z(n216) );
  INV_X1 U249 ( .A(n3998), .ZN(n3995) );
  INV_X4 U251 ( .A(n3825), .ZN(n59) );
  NAND2_X1 U252 ( .A1(n514), .A2(n516), .ZN(n1185) );
  INV_X2 U253 ( .A(n2269), .ZN(n2091) );
  INV_X2 U256 ( .A(n1989), .ZN(n60) );
  XNOR2_X1 U257 ( .A(n3756), .B(n3757), .ZN(n3759) );
  INV_X2 U258 ( .A(n4024), .ZN(n61) );
  NAND2_X2 U259 ( .A1(n1530), .A2(n1529), .ZN(n3736) );
  INV_X2 U260 ( .A(n3817), .ZN(n3813) );
  INV_X4 U261 ( .A(n3753), .ZN(n62) );
  INV_X2 U262 ( .A(n3685), .ZN(n3686) );
  INV_X2 U263 ( .A(n3610), .ZN(n1848) );
  NOR2_X2 U265 ( .A1(n3099), .A2(n3098), .ZN(n3561) );
  INV_X2 U266 ( .A(n2676), .ZN(n850) );
  INV_X2 U267 ( .A(n684), .ZN(n3230) );
  INV_X4 U268 ( .A(n2652), .ZN(n63) );
  INV_X2 U269 ( .A(n2148), .ZN(n1579) );
  NOR2_X2 U270 ( .A1(n1973), .A2(n3766), .ZN(n1970) );
  INV_X2 U272 ( .A(n2326), .ZN(n2008) );
  INV_X2 U274 ( .A(n3374), .ZN(n3376) );
  INV_X4 U276 ( .A(n3173), .ZN(n64) );
  INV_X2 U278 ( .A(n942), .ZN(n782) );
  NAND2_X2 U279 ( .A1(n1378), .A2(n1643), .ZN(n824) );
  INV_X2 U280 ( .A(n2992), .ZN(n65) );
  NAND2_X2 U282 ( .A1(n2330), .A2(n3256), .ZN(n1365) );
  INV_X4 U283 ( .A(n1644), .ZN(n66) );
  INV_X4 U285 ( .A(n1222), .ZN(n68) );
  INV_X2 U286 ( .A(n2770), .ZN(n2769) );
  INV_X2 U287 ( .A(n2599), .ZN(n732) );
  INV_X4 U288 ( .A(n366), .ZN(n69) );
  OR2_X2 U291 ( .A1(n3355), .A2(n1777), .ZN(n471) );
  INV_X2 U292 ( .A(n709), .ZN(n3048) );
  INV_X2 U293 ( .A(n2745), .ZN(n2747) );
  INV_X4 U295 ( .A(n3442), .ZN(n70) );
  INV_X2 U296 ( .A(n3400), .ZN(n1560) );
  NOR2_X2 U297 ( .A1(n3346), .A2(n3345), .ZN(n3365) );
  NAND2_X2 U298 ( .A1(n3346), .A2(n3345), .ZN(n3363) );
  INV_X4 U299 ( .A(n2966), .ZN(n71) );
  INV_X2 U300 ( .A(n2493), .ZN(n2490) );
  BUF_X4 U301 ( .A(n3555), .Z(n1666) );
  INV_X2 U302 ( .A(n1680), .ZN(n574) );
  INV_X4 U303 ( .A(n2973), .ZN(n72) );
  INV_X2 U304 ( .A(n412), .ZN(n413) );
  INV_X2 U308 ( .A(n2532), .ZN(n1376) );
  INV_X4 U309 ( .A(n1686), .ZN(n73) );
  INV_X2 U311 ( .A(n2626), .ZN(n2628) );
  XNOR2_X1 U312 ( .A(n3486), .B(n3485), .ZN(n3488) );
  INV_X2 U313 ( .A(n2624), .ZN(n2623) );
  NAND2_X2 U314 ( .A1(n262), .A2(n263), .ZN(n687) );
  INV_X2 U315 ( .A(n1739), .ZN(n1592) );
  INV_X2 U316 ( .A(n2137), .ZN(n1331) );
  INV_X2 U319 ( .A(n2404), .ZN(n604) );
  NAND2_X1 U320 ( .A1(n1547), .A2(n1548), .ZN(n1550) );
  INV_X2 U321 ( .A(n2511), .ZN(n1332) );
  NOR2_X1 U322 ( .A1(n2718), .A2(n2717), .ZN(n2723) );
  NAND2_X1 U323 ( .A1(n2339), .A2(n2302), .ZN(n127) );
  INV_X2 U325 ( .A(n261), .ZN(n262) );
  INV_X2 U327 ( .A(n3347), .ZN(n3350) );
  INV_X2 U329 ( .A(n3191), .ZN(n3195) );
  AND2_X2 U332 ( .A1(n3404), .A2(n1692), .ZN(n461) );
  INV_X2 U335 ( .A(n2510), .ZN(n1333) );
  AND2_X1 U336 ( .A1(n3545), .A2(n3543), .ZN(n464) );
  INV_X2 U338 ( .A(n1397), .ZN(n1277) );
  AND2_X2 U339 ( .A1(n3251), .A2(n3250), .ZN(n447) );
  OAI21_X1 U340 ( .B1(n1106), .B2(n1105), .A(n2546), .ZN(n1104) );
  NAND2_X2 U341 ( .A1(n583), .A2(n582), .ZN(n2523) );
  INV_X2 U342 ( .A(n3418), .ZN(n1552) );
  INV_X2 U343 ( .A(n1768), .ZN(n1767) );
  NOR2_X2 U344 ( .A1(n2664), .A2(n2616), .ZN(n1286) );
  INV_X4 U346 ( .A(n2722), .ZN(n75) );
  INV_X2 U347 ( .A(n3246), .ZN(n1634) );
  NAND2_X2 U348 ( .A1(n2265), .A2(n2266), .ZN(n645) );
  INV_X4 U349 ( .A(n2993), .ZN(n76) );
  INV_X2 U350 ( .A(n2990), .ZN(n1454) );
  INV_X2 U352 ( .A(n4178), .ZN(n77) );
  OR2_X2 U353 ( .A1(n2707), .A2(n2706), .ZN(n2711) );
  INV_X2 U356 ( .A(n2790), .ZN(n2784) );
  NAND2_X2 U357 ( .A1(n3391), .A2(n3390), .ZN(n3418) );
  NAND2_X1 U360 ( .A1(n2130), .A2(n2988), .ZN(n2888) );
  AND2_X1 U361 ( .A1(n2753), .A2(n2714), .ZN(n2693) );
  NOR2_X2 U362 ( .A1(n460), .A2(n2424), .ZN(n2428) );
  NAND2_X2 U363 ( .A1(n2410), .A2(n4055), .ZN(n2510) );
  INV_X2 U365 ( .A(n2202), .ZN(n1308) );
  INV_X2 U366 ( .A(n2513), .ZN(n78) );
  INV_X2 U367 ( .A(n2753), .ZN(n2701) );
  NAND2_X1 U369 ( .A1(n487), .A2(n4041), .ZN(n2896) );
  INV_X2 U370 ( .A(n2455), .ZN(n2456) );
  INV_X2 U371 ( .A(n2956), .ZN(n1015) );
  NAND2_X2 U373 ( .A1(n2681), .A2(n2680), .ZN(n3595) );
  NAND2_X1 U374 ( .A1(n2793), .A2(n2270), .ZN(n2794) );
  INV_X2 U375 ( .A(n2408), .ZN(n2410) );
  INV_X2 U376 ( .A(n733), .ZN(n603) );
  NAND2_X2 U378 ( .A1(n2660), .A2(n2659), .ZN(n2757) );
  INV_X2 U381 ( .A(n2546), .ZN(n80) );
  INV_X4 U382 ( .A(n150), .ZN(n2201) );
  INV_X4 U383 ( .A(n3467), .ZN(n81) );
  INV_X2 U384 ( .A(n622), .ZN(n3079) );
  NAND3_X1 U385 ( .A1(n2807), .A2(n3202), .A3(n2806), .ZN(n2808) );
  NAND2_X1 U386 ( .A1(n230), .A2(n1784), .ZN(n228) );
  INV_X2 U387 ( .A(n2478), .ZN(n82) );
  NOR2_X1 U388 ( .A1(n327), .A2(n326), .ZN(n325) );
  INV_X4 U389 ( .A(n2022), .ZN(n2736) );
  INV_X1 U390 ( .A(n3500), .ZN(n3527) );
  INV_X4 U391 ( .A(n3051), .ZN(n83) );
  AND2_X2 U392 ( .A1(n2221), .A2(n2222), .ZN(n469) );
  AND2_X2 U393 ( .A1(n560), .A2(n2809), .ZN(n443) );
  INV_X4 U395 ( .A(n241), .ZN(n2296) );
  MUX2_X1 U397 ( .A(n3839), .B(n3113), .S(a[24]), .Z(n3639) );
  INV_X4 U399 ( .A(n1720), .ZN(n1721) );
  INV_X2 U403 ( .A(n3077), .ZN(n2094) );
  OR2_X2 U406 ( .A1(n1370), .A2(n3217), .ZN(n453) );
  NAND2_X1 U407 ( .A1(n2787), .A2(n2217), .ZN(n2216) );
  INV_X8 U408 ( .A(n3310), .ZN(n85) );
  INV_X8 U410 ( .A(n2084), .ZN(n86) );
  AND2_X1 U411 ( .A1(n1890), .A2(a[9]), .ZN(n474) );
  INV_X8 U412 ( .A(n3200), .ZN(n87) );
  AND2_X2 U414 ( .A1(n2803), .A2(n2802), .ZN(n1056) );
  AND2_X2 U415 ( .A1(n3067), .A2(n2825), .ZN(n2390) );
  INV_X2 U416 ( .A(n2411), .ZN(n1231) );
  INV_X4 U418 ( .A(n2941), .ZN(n88) );
  AND2_X2 U421 ( .A1(n2982), .A2(n3124), .ZN(n427) );
  AND2_X2 U422 ( .A1(n3065), .A2(n3139), .ZN(n187) );
  AND2_X2 U423 ( .A1(n2982), .A2(a[21]), .ZN(n463) );
  NAND2_X2 U424 ( .A1(n99), .A2(b[14]), .ZN(n2824) );
  NOR2_X2 U427 ( .A1(n3468), .A2(n2907), .ZN(n2908) );
  NAND2_X2 U429 ( .A1(n291), .A2(n2785), .ZN(n1024) );
  INV_X4 U431 ( .A(n2356), .ZN(n95) );
  INV_X2 U432 ( .A(n2438), .ZN(n96) );
  INV_X2 U435 ( .A(n2407), .ZN(n98) );
  INV_X4 U436 ( .A(n1784), .ZN(n99) );
  INV_X4 U437 ( .A(a[2]), .ZN(n2355) );
  INV_X4 U438 ( .A(n3468), .ZN(n100) );
  NAND2_X2 U439 ( .A1(n414), .A2(n413), .ZN(n115) );
  NAND3_X2 U440 ( .A1(n3111), .A2(n667), .A3(n3110), .ZN(n414) );
  INV_X4 U441 ( .A(n2853), .ZN(n504) );
  NAND2_X2 U442 ( .A1(n1220), .A2(n1796), .ZN(n2173) );
  NAND2_X2 U443 ( .A1(n3382), .A2(n612), .ZN(n1220) );
  NAND2_X2 U444 ( .A1(n831), .A2(n99), .ZN(n1063) );
  INV_X4 U445 ( .A(n2830), .ZN(n1720) );
  NOR2_X2 U446 ( .A1(n3094), .A2(n1222), .ZN(n1708) );
  INV_X4 U447 ( .A(n3093), .ZN(n3094) );
  NAND2_X2 U448 ( .A1(n1066), .A2(n1065), .ZN(n3093) );
  NAND2_X2 U449 ( .A1(n101), .A2(n1506), .ZN(n2286) );
  NAND2_X2 U450 ( .A1(n1505), .A2(n2971), .ZN(n101) );
  NOR2_X2 U452 ( .A1(n89), .A2(n2899), .ZN(n877) );
  AOI22_X2 U453 ( .A1(n1217), .A2(n3203), .B1(n3080), .B2(n58), .ZN(n2899) );
  NAND2_X2 U455 ( .A1(n102), .A2(n3556), .ZN(n2238) );
  NAND2_X2 U460 ( .A1(n1729), .A2(n3051), .ZN(n1728) );
  NOR2_X4 U463 ( .A1(n1265), .A2(n2385), .ZN(n3044) );
  NAND2_X2 U464 ( .A1(n104), .A2(n2865), .ZN(n2869) );
  NAND2_X2 U465 ( .A1(n4058), .A2(n914), .ZN(n104) );
  BUF_X4 U466 ( .A(n241), .Z(n105) );
  NAND2_X2 U468 ( .A1(n107), .A2(n1454), .ZN(n489) );
  INV_X2 U469 ( .A(n2040), .ZN(n107) );
  NAND2_X2 U470 ( .A1(n876), .A2(n875), .ZN(n2040) );
  INV_X4 U471 ( .A(n571), .ZN(n3644) );
  INV_X4 U473 ( .A(n3893), .ZN(n3898) );
  OAI21_X2 U474 ( .B1(n211), .B2(n210), .A(n2950), .ZN(n3173) );
  OAI21_X2 U476 ( .B1(n751), .B2(n1299), .A(n3175), .ZN(n3570) );
  NOR2_X2 U480 ( .A1(n1161), .A2(n2943), .ZN(n2185) );
  NAND2_X2 U481 ( .A1(n1213), .A2(n1212), .ZN(n1161) );
  NAND2_X2 U482 ( .A1(n109), .A2(n4071), .ZN(n1904) );
  NAND2_X2 U484 ( .A1(n3571), .A2(n3570), .ZN(n3911) );
  NAND2_X2 U485 ( .A1(n2054), .A2(n2055), .ZN(n1498) );
  INV_X2 U486 ( .A(n3134), .ZN(n1210) );
  NAND2_X2 U487 ( .A1(n1046), .A2(n1045), .ZN(n3134) );
  INV_X4 U488 ( .A(n3228), .ZN(n1036) );
  NAND2_X2 U489 ( .A1(n110), .A2(n3095), .ZN(n1502) );
  INV_X4 U491 ( .A(n661), .ZN(n1620) );
  NAND2_X1 U492 ( .A1(n105), .A2(n3202), .ZN(n2436) );
  NAND2_X2 U493 ( .A1(n111), .A2(a[25]), .ZN(n2614) );
  NAND2_X2 U495 ( .A1(n111), .A2(a[17]), .ZN(n1948) );
  NAND2_X2 U496 ( .A1(n111), .A2(n2356), .ZN(n2183) );
  NAND2_X1 U497 ( .A1(n2070), .A2(a[1]), .ZN(n3425) );
  NAND2_X2 U498 ( .A1(n3124), .A2(n111), .ZN(n799) );
  NAND2_X2 U499 ( .A1(n111), .A2(a[7]), .ZN(n1732) );
  NAND2_X1 U500 ( .A1(n111), .A2(n1784), .ZN(n301) );
  NAND2_X1 U502 ( .A1(n1784), .A2(n111), .ZN(n1064) );
  NAND2_X2 U503 ( .A1(n56), .A2(n111), .ZN(n834) );
  NAND2_X2 U504 ( .A1(n111), .A2(a[24]), .ZN(n895) );
  INV_X8 U505 ( .A(n3206), .ZN(n111) );
  NAND2_X4 U508 ( .A1(n1342), .A2(n115), .ZN(n1223) );
  NOR2_X2 U509 ( .A1(n116), .A2(n2374), .ZN(n2377) );
  BUF_X4 U510 ( .A(n1834), .Z(n117) );
  INV_X4 U511 ( .A(n1834), .ZN(n2654) );
  NAND2_X2 U512 ( .A1(n241), .A2(n1834), .ZN(n571) );
  NAND2_X4 U513 ( .A1(n249), .A2(n2924), .ZN(n1834) );
  NAND2_X2 U514 ( .A1(n822), .A2(n821), .ZN(n3337) );
  NAND2_X2 U515 ( .A1(n824), .A2(n823), .ZN(n3338) );
  NAND4_X1 U516 ( .A1(n824), .A2(n4140), .A3(n821), .A4(n823), .ZN(n612) );
  NAND2_X2 U517 ( .A1(n1101), .A2(n3347), .ZN(n821) );
  NAND2_X2 U519 ( .A1(n3354), .A2(n624), .ZN(n823) );
  NAND2_X2 U520 ( .A1(n1160), .A2(n817), .ZN(n436) );
  NAND2_X2 U521 ( .A1(n123), .A2(n121), .ZN(n817) );
  INV_X2 U523 ( .A(n121), .ZN(n118) );
  INV_X2 U524 ( .A(n123), .ZN(n119) );
  OAI22_X2 U526 ( .A1(n916), .A2(n3204), .B1(n3538), .B2(n1303), .ZN(n124) );
  AOI21_X2 U527 ( .B1(n4040), .B2(n1100), .A(n1099), .ZN(n121) );
  AOI21_X2 U528 ( .B1(n825), .B2(n826), .A(n124), .ZN(n123) );
  NOR2_X2 U530 ( .A1(n127), .A2(n1558), .ZN(n1557) );
  NAND2_X4 U534 ( .A1(n130), .A2(n128), .ZN(n1686) );
  NAND2_X2 U537 ( .A1(n1688), .A2(n2435), .ZN(n2513) );
  NAND2_X2 U538 ( .A1(n2512), .A2(n131), .ZN(n130) );
  NAND3_X1 U539 ( .A1(n1688), .A2(n2435), .A3(n1687), .ZN(n131) );
  NAND3_X2 U540 ( .A1(n1689), .A2(n2023), .A3(n4053), .ZN(n2512) );
  NAND2_X2 U542 ( .A1(n1558), .A2(n2514), .ZN(n133) );
  NAND2_X4 U544 ( .A1(n2002), .A2(n2001), .ZN(n3933) );
  OAI21_X2 U545 ( .B1(n135), .B2(n2528), .A(n134), .ZN(n2001) );
  NAND2_X1 U546 ( .A1(n743), .A2(n1893), .ZN(n134) );
  NOR2_X1 U547 ( .A1(n743), .A2(n1893), .ZN(n135) );
  NAND2_X2 U548 ( .A1(n137), .A2(n136), .ZN(n2002) );
  NAND3_X1 U549 ( .A1(n1372), .A2(n2606), .A3(n1373), .ZN(n136) );
  NAND2_X2 U550 ( .A1(n1133), .A2(n1134), .ZN(n137) );
  NOR2_X4 U551 ( .A1(n1990), .A2(n2191), .ZN(n931) );
  NAND2_X4 U552 ( .A1(n139), .A2(n138), .ZN(n2191) );
  INV_X2 U553 ( .A(n933), .ZN(n138) );
  NAND2_X2 U554 ( .A1(n141), .A2(n140), .ZN(n1990) );
  NAND3_X1 U555 ( .A1(n1356), .A2(n2528), .A3(n1355), .ZN(n140) );
  NAND2_X2 U556 ( .A1(n764), .A2(n744), .ZN(n141) );
  NAND3_X2 U557 ( .A1(n3674), .A2(n3673), .A3(n3672), .ZN(\d[38]_BAR ) );
  INV_X2 U559 ( .A(n1876), .ZN(n2043) );
  NAND2_X2 U560 ( .A1(n4181), .A2(n142), .ZN(n1876) );
  NOR2_X2 U561 ( .A1(n2922), .A2(n4182), .ZN(n1961) );
  NOR2_X2 U562 ( .A1(n143), .A2(n142), .ZN(n2039) );
  AOI22_X2 U563 ( .A1(n2818), .A2(n2817), .B1(n2816), .B2(n1537), .ZN(n142) );
  NAND2_X2 U564 ( .A1(n2135), .A2(n2134), .ZN(n143) );
  OAI21_X2 U565 ( .B1(n2877), .B2(n201), .A(n626), .ZN(n2922) );
  NAND2_X2 U566 ( .A1(n527), .A2(n2875), .ZN(n626) );
  NAND2_X2 U567 ( .A1(n1877), .A2(n1876), .ZN(n144) );
  INV_X2 U568 ( .A(n2922), .ZN(n145) );
  NAND2_X2 U569 ( .A1(n146), .A2(n2397), .ZN(n1656) );
  NAND2_X2 U570 ( .A1(n2398), .A2(n146), .ZN(n3633) );
  NAND2_X2 U571 ( .A1(n3662), .A2(n146), .ZN(n3673) );
  INV_X4 U572 ( .A(n3863), .ZN(n146) );
  NOR2_X1 U573 ( .A1(n147), .A2(n3602), .ZN(n3626) );
  NAND3_X2 U574 ( .A1(n147), .A2(n3929), .A3(n3928), .ZN(n3930) );
  INV_X4 U576 ( .A(n2852), .ZN(n2903) );
  NAND3_X2 U578 ( .A1(n1173), .A2(n1569), .A3(n1174), .ZN(n970) );
  NAND2_X2 U581 ( .A1(n2012), .A2(n1578), .ZN(n818) );
  NAND3_X2 U582 ( .A1(n828), .A2(n1607), .A3(n1606), .ZN(n2012) );
  NAND2_X2 U583 ( .A1(n870), .A2(n148), .ZN(n588) );
  NAND3_X2 U584 ( .A1(n490), .A2(n1486), .A3(n3025), .ZN(n148) );
  NAND2_X2 U585 ( .A1(n493), .A2(n494), .ZN(n492) );
  INV_X2 U586 ( .A(n1230), .ZN(n2960) );
  NAND2_X2 U588 ( .A1(n2031), .A2(n2082), .ZN(n2037) );
  INV_X2 U589 ( .A(n1449), .ZN(n150) );
  INV_X2 U590 ( .A(n1914), .ZN(n2894) );
  NAND2_X2 U593 ( .A1(n1918), .A2(n20), .ZN(n151) );
  NAND2_X2 U594 ( .A1(n152), .A2(n3169), .ZN(n3226) );
  NAND3_X2 U595 ( .A1(n1304), .A2(n2036), .A3(n2037), .ZN(n152) );
  NAND2_X2 U596 ( .A1(n3606), .A2(n1636), .ZN(n1737) );
  NAND3_X2 U597 ( .A1(n1637), .A2(n3569), .A3(n4004), .ZN(n3606) );
  NOR2_X2 U601 ( .A1(n276), .A2(n2945), .ZN(n275) );
  NAND2_X2 U602 ( .A1(n217), .A2(n1684), .ZN(n276) );
  BUF_X4 U603 ( .A(n86), .Z(n155) );
  NOR2_X4 U604 ( .A1(n156), .A2(n3027), .ZN(n1131) );
  NAND2_X1 U610 ( .A1(n3328), .A2(n3118), .ZN(n2349) );
  NAND2_X2 U611 ( .A1(n3453), .A2(a[19]), .ZN(n555) );
  NOR2_X2 U612 ( .A1(n22), .A2(n1623), .ZN(n1622) );
  INV_X8 U613 ( .A(n1913), .ZN(n1227) );
  INV_X4 U614 ( .A(n158), .ZN(n1399) );
  NOR2_X2 U615 ( .A1(n1944), .A2(n2995), .ZN(n158) );
  NAND3_X2 U616 ( .A1(n2299), .A2(n1081), .A3(n2228), .ZN(n1317) );
  NOR2_X2 U618 ( .A1(n3333), .A2(n3332), .ZN(n159) );
  AOI21_X2 U619 ( .B1(n3333), .B2(n3332), .A(n3334), .ZN(n160) );
  NAND2_X2 U620 ( .A1(n2769), .A2(n1452), .ZN(n2773) );
  NAND2_X2 U621 ( .A1(n1411), .A2(n3377), .ZN(n1413) );
  AOI22_X2 U623 ( .A1(n3921), .A2(n3920), .B1(n3919), .B2(n3918), .ZN(n3922)
         );
  NAND2_X2 U624 ( .A1(n161), .A2(n2319), .ZN(n188) );
  NAND2_X2 U629 ( .A1(n1616), .A2(n1615), .ZN(n611) );
  NOR2_X2 U630 ( .A1(n1286), .A2(n2106), .ZN(n1855) );
  OAI21_X2 U633 ( .B1(n162), .B2(n1627), .A(n1626), .ZN(n808) );
  NAND2_X2 U634 ( .A1(n1956), .A2(n1957), .ZN(n162) );
  NOR2_X4 U635 ( .A1(n771), .A2(n3296), .ZN(n2279) );
  AOI22_X2 U636 ( .A1(n3190), .A2(n3189), .B1(n1282), .B2(n3188), .ZN(n3197)
         );
  NAND3_X2 U637 ( .A1(n175), .A2(n3738), .A3(n3911), .ZN(n1509) );
  NOR2_X2 U638 ( .A1(n2329), .A2(n3298), .ZN(n220) );
  NOR2_X2 U640 ( .A1(n163), .A2(n259), .ZN(n258) );
  NAND2_X4 U642 ( .A1(n385), .A2(n3282), .ZN(n3290) );
  NOR3_X2 U643 ( .A1(n665), .A2(n663), .A3(n664), .ZN(n2319) );
  NAND2_X2 U645 ( .A1(n2995), .A2(n1944), .ZN(n1398) );
  NAND2_X2 U646 ( .A1(n1258), .A2(n1259), .ZN(n1944) );
  NAND3_X2 U647 ( .A1(n4210), .A2(n4069), .A3(n746), .ZN(n2528) );
  XNOR2_X2 U648 ( .A(n164), .B(n3370), .ZN(n3806) );
  AOI22_X2 U649 ( .A1(n867), .A2(n66), .B1(n1644), .B2(n3559), .ZN(n164) );
  AOI22_X2 U650 ( .A1(n2263), .A2(n1661), .B1(n1711), .B2(n509), .ZN(n1589) );
  INV_X4 U651 ( .A(n2906), .ZN(n3409) );
  NAND2_X4 U652 ( .A1(n2128), .A2(n3290), .ZN(n2127) );
  NAND3_X2 U653 ( .A1(n165), .A2(n965), .A3(n964), .ZN(n963) );
  INV_X2 U654 ( .A(n967), .ZN(n165) );
  NAND2_X2 U655 ( .A1(n1562), .A2(n1561), .ZN(n967) );
  NOR2_X4 U658 ( .A1(n570), .A2(n166), .ZN(n3340) );
  NAND2_X2 U659 ( .A1(n568), .A2(n569), .ZN(n166) );
  NAND2_X2 U660 ( .A1(n167), .A2(n1415), .ZN(n1833) );
  NAND2_X2 U661 ( .A1(n1097), .A2(n1414), .ZN(n167) );
  NOR2_X4 U662 ( .A1(n168), .A2(n3393), .ZN(n3435) );
  NAND2_X2 U663 ( .A1(n2184), .A2(n2183), .ZN(n168) );
  NAND2_X2 U664 ( .A1(n831), .A2(n3407), .ZN(n1731) );
  OAI21_X2 U665 ( .B1(n3305), .B2(n3304), .A(n2366), .ZN(n2363) );
  AOI21_X2 U666 ( .B1(n1290), .B2(n3062), .A(n3059), .ZN(n1382) );
  NOR2_X2 U667 ( .A1(n3797), .A2(n3810), .ZN(n3819) );
  AOI21_X2 U668 ( .B1(n3028), .B2(n3029), .A(n3030), .ZN(n3039) );
  AOI22_X2 U669 ( .A1(n689), .A2(n2982), .B1(n3016), .B2(n1088), .ZN(n3030) );
  NOR2_X2 U670 ( .A1(n3793), .A2(n3792), .ZN(n3829) );
  NAND2_X2 U671 ( .A1(n1438), .A2(n1437), .ZN(n3793) );
  INV_X2 U673 ( .A(n508), .ZN(n169) );
  NAND2_X2 U674 ( .A1(n510), .A2(n509), .ZN(n508) );
  NAND2_X4 U676 ( .A1(n827), .A2(n4179), .ZN(n509) );
  NAND2_X4 U677 ( .A1(n538), .A2(n509), .ZN(n2263) );
  NAND2_X2 U678 ( .A1(n1124), .A2(n3089), .ZN(n1864) );
  AOI22_X2 U679 ( .A1(n2113), .A2(n219), .B1(n266), .B2(n19), .ZN(n2285) );
  NAND2_X2 U680 ( .A1(n1460), .A2(n1461), .ZN(n1074) );
  NAND2_X1 U682 ( .A1(n2306), .A2(n1804), .ZN(n3731) );
  NOR2_X2 U683 ( .A1(n2308), .A2(n2307), .ZN(n2306) );
  NOR2_X1 U685 ( .A1(n1558), .A2(n2518), .ZN(n2515) );
  NAND3_X2 U686 ( .A1(n1004), .A2(n171), .A3(n170), .ZN(n1003) );
  NAND2_X2 U688 ( .A1(n333), .A2(n1005), .ZN(n171) );
  NOR2_X2 U689 ( .A1(n3906), .A2(n62), .ZN(n466) );
  NAND2_X2 U692 ( .A1(n1174), .A2(n1173), .ZN(n620) );
  NAND2_X2 U693 ( .A1(n621), .A2(n71), .ZN(n1174) );
  AOI21_X2 U694 ( .B1(n2473), .B2(n2474), .A(n35), .ZN(n1159) );
  NAND2_X2 U695 ( .A1(n4025), .A2(n4019), .ZN(n3699) );
  NOR2_X2 U697 ( .A1(n1102), .A2(n3291), .ZN(n369) );
  NAND2_X2 U698 ( .A1(n372), .A2(n373), .ZN(n1102) );
  INV_X4 U699 ( .A(n2504), .ZN(n2253) );
  NAND2_X2 U701 ( .A1(n2653), .A2(n728), .ZN(n727) );
  NAND3_X2 U702 ( .A1(n731), .A2(n732), .A3(n1496), .ZN(n2653) );
  NAND3_X2 U705 ( .A1(n2465), .A2(n174), .A3(n173), .ZN(n2469) );
  NAND3_X2 U707 ( .A1(n954), .A2(n2105), .A3(n2013), .ZN(n630) );
  NAND2_X4 U710 ( .A1(n2127), .A2(n1539), .ZN(n1483) );
  INV_X2 U711 ( .A(n384), .ZN(n175) );
  INV_X1 U712 ( .A(n675), .ZN(n260) );
  NAND2_X4 U713 ( .A1(n388), .A2(n389), .ZN(n3258) );
  NAND2_X2 U714 ( .A1(n2697), .A2(n3431), .ZN(n1179) );
  NAND2_X2 U715 ( .A1(n176), .A2(n3252), .ZN(n389) );
  INV_X2 U716 ( .A(n1367), .ZN(n176) );
  NAND3_X2 U717 ( .A1(n1179), .A2(n1175), .A3(n1176), .ZN(n1367) );
  NAND2_X2 U718 ( .A1(n177), .A2(n1512), .ZN(n3353) );
  NOR2_X2 U722 ( .A1(n3791), .A2(n2269), .ZN(n3887) );
  NOR2_X2 U723 ( .A1(n3810), .A2(n2089), .ZN(n3791) );
  NOR2_X4 U726 ( .A1(n3412), .A2(n178), .ZN(n721) );
  NAND2_X2 U728 ( .A1(n1209), .A2(n1221), .ZN(n179) );
  INV_X1 U731 ( .A(n4021), .ZN(n181) );
  NOR2_X2 U732 ( .A1(n3730), .A2(n3693), .ZN(n2397) );
  NAND3_X2 U734 ( .A1(n1166), .A2(n2789), .A3(n469), .ZN(n802) );
  NAND2_X2 U735 ( .A1(n182), .A2(n3882), .ZN(\d[39] ) );
  OAI22_X2 U736 ( .A1(n3862), .A2(n302), .B1(n3861), .B2(n3860), .ZN(n182) );
  INV_X4 U737 ( .A(n432), .ZN(n560) );
  NOR2_X2 U741 ( .A1(n3713), .A2(n3863), .ZN(n3727) );
  XNOR2_X2 U744 ( .A(n3339), .B(n991), .ZN(n1964) );
  NAND2_X2 U745 ( .A1(n993), .A2(n992), .ZN(n3339) );
  OAI21_X2 U746 ( .B1(n3275), .B2(n2392), .A(n184), .ZN(n3287) );
  INV_X2 U747 ( .A(n3274), .ZN(n184) );
  NOR2_X2 U748 ( .A1(n1696), .A2(n3242), .ZN(n3274) );
  OAI22_X2 U749 ( .A1(n2084), .A2(n3534), .B1(n3328), .B2(a[3]), .ZN(n994) );
  BUF_X4 U750 ( .A(n3777), .Z(n185) );
  NAND3_X2 U751 ( .A1(n3072), .A2(n3071), .A3(n186), .ZN(n622) );
  NAND3_X1 U752 ( .A1(n3070), .A2(n187), .A3(n2193), .ZN(n186) );
  NAND2_X2 U753 ( .A1(n894), .A2(n3340), .ZN(n1473) );
  NAND3_X2 U754 ( .A1(n188), .A2(n3785), .A3(n3799), .ZN(n1260) );
  NAND2_X2 U756 ( .A1(n366), .A2(n2564), .ZN(n189) );
  AOI21_X2 U757 ( .B1(n1243), .B2(n3754), .A(n1479), .ZN(n3755) );
  NOR2_X2 U758 ( .A1(n827), .A2(n3090), .ZN(n539) );
  NAND2_X4 U759 ( .A1(n917), .A2(n3088), .ZN(n827) );
  INV_X4 U760 ( .A(n1323), .ZN(n559) );
  AOI21_X2 U761 ( .B1(n2992), .B2(n2976), .A(n2975), .ZN(n2046) );
  NAND2_X2 U762 ( .A1(n903), .A2(n900), .ZN(n2976) );
  NAND2_X2 U764 ( .A1(n191), .A2(n206), .ZN(n1638) );
  NAND2_X2 U765 ( .A1(n1226), .A2(n3565), .ZN(n191) );
  NAND2_X2 U766 ( .A1(n596), .A2(n967), .ZN(n1691) );
  NOR2_X2 U768 ( .A1(n1181), .A2(n458), .ZN(n1688) );
  NOR2_X1 U769 ( .A1(n3026), .A2(n2913), .ZN(n2914) );
  NAND2_X2 U770 ( .A1(n262), .A2(n2544), .ZN(n367) );
  INV_X2 U771 ( .A(n1316), .ZN(n435) );
  NAND2_X2 U772 ( .A1(n193), .A2(n192), .ZN(n1316) );
  INV_X2 U773 ( .A(n1363), .ZN(n192) );
  INV_X2 U774 ( .A(n3605), .ZN(n193) );
  AOI21_X2 U775 ( .B1(n3730), .B2(n3704), .A(n3703), .ZN(n3705) );
  INV_X4 U776 ( .A(n3572), .ZN(n332) );
  NAND2_X4 U779 ( .A1(n3966), .A2(n3299), .ZN(n331) );
  INV_X8 U780 ( .A(n331), .ZN(n4018) );
  NAND2_X2 U781 ( .A1(n3200), .A2(n2407), .ZN(n556) );
  NOR2_X4 U784 ( .A1(n3730), .A2(n2060), .ZN(n2396) );
  NAND2_X2 U785 ( .A1(n196), .A2(n3197), .ZN(n2041) );
  NAND3_X2 U786 ( .A1(n3195), .A2(n3196), .A3(n3192), .ZN(n196) );
  NOR2_X2 U787 ( .A1(n197), .A2(n2942), .ZN(n3159) );
  OAI21_X2 U789 ( .B1(n2964), .B2(n2965), .A(n198), .ZN(n3106) );
  NAND2_X1 U792 ( .A1(n1227), .A2(n1340), .ZN(n2225) );
  NAND2_X2 U793 ( .A1(n199), .A2(n3108), .ZN(n1741) );
  NAND3_X2 U794 ( .A1(n1742), .A2(n1007), .A3(n1008), .ZN(n199) );
  NAND2_X2 U795 ( .A1(n200), .A2(n1052), .ZN(n1051) );
  NAND2_X2 U796 ( .A1(n1054), .A2(n1053), .ZN(n200) );
  INV_X4 U797 ( .A(n748), .ZN(n3070) );
  XOR2_X2 U798 ( .A(n3498), .B(a[11]), .Z(n3007) );
  NOR2_X4 U799 ( .A1(n3909), .A2(n3911), .ZN(n661) );
  NAND2_X4 U801 ( .A1(n1596), .A2(n1597), .ZN(n1599) );
  NAND2_X2 U802 ( .A1(n656), .A2(n655), .ZN(n654) );
  NAND2_X2 U803 ( .A1(n705), .A2(n64), .ZN(n656) );
  NAND2_X2 U804 ( .A1(n3854), .A2(n3924), .ZN(n3602) );
  XNOR2_X2 U806 ( .A(n2499), .B(n2620), .ZN(n2600) );
  NAND2_X2 U807 ( .A1(n204), .A2(n203), .ZN(n2497) );
  NAND2_X2 U808 ( .A1(a[17]), .A2(n2022), .ZN(n203) );
  NAND2_X2 U811 ( .A1(n1964), .A2(n1963), .ZN(n1472) );
  NOR2_X2 U812 ( .A1(n599), .A2(n3817), .ZN(n819) );
  OAI21_X2 U813 ( .B1(n2196), .B2(n3787), .A(n2194), .ZN(n599) );
  BUF_X4 U814 ( .A(n3468), .Z(n205) );
  NAND2_X2 U816 ( .A1(n3239), .A2(n3238), .ZN(n1517) );
  INV_X2 U817 ( .A(n3566), .ZN(n206) );
  OAI21_X2 U818 ( .B1(n2007), .B2(n3564), .A(n3567), .ZN(n3566) );
  NAND2_X2 U820 ( .A1(n4037), .A2(n911), .ZN(n207) );
  NAND2_X2 U821 ( .A1(n1844), .A2(n3084), .ZN(n3361) );
  NAND2_X2 U822 ( .A1(n1424), .A2(n1423), .ZN(n1844) );
  NAND3_X2 U823 ( .A1(n551), .A2(n552), .A3(n250), .ZN(n550) );
  NAND2_X2 U824 ( .A1(n2984), .A2(n2985), .ZN(n1457) );
  NAND2_X2 U825 ( .A1(n3052), .A2(n3051), .ZN(n1425) );
  NAND3_X2 U827 ( .A1(n1459), .A2(n1575), .A3(n1574), .ZN(n1461) );
  NAND2_X2 U829 ( .A1(n2117), .A2(n1418), .ZN(n1707) );
  NAND2_X2 U830 ( .A1(n1609), .A2(n1608), .ZN(n1418) );
  OAI21_X2 U831 ( .B1(n1937), .B2(n2297), .A(n3102), .ZN(n2117) );
  NOR2_X2 U833 ( .A1(n209), .A2(n4152), .ZN(n1758) );
  NOR2_X2 U834 ( .A1(n1830), .A2(n3022), .ZN(n209) );
  OAI21_X2 U835 ( .B1(n302), .B2(n239), .A(n3657), .ZN(n3674) );
  NOR2_X2 U836 ( .A1(n977), .A2(n2948), .ZN(n210) );
  INV_X2 U837 ( .A(n2949), .ZN(n211) );
  NAND2_X2 U838 ( .A1(n3945), .A2(n3946), .ZN(n3948) );
  INV_X4 U840 ( .A(n212), .ZN(n1607) );
  NOR2_X2 U841 ( .A1(n726), .A2(n1589), .ZN(n212) );
  NOR2_X4 U842 ( .A1(n332), .A2(n661), .ZN(n3966) );
  INV_X4 U843 ( .A(b[11]), .ZN(n1315) );
  NOR2_X4 U844 ( .A1(n3129), .A2(n3125), .ZN(n1261) );
  NAND2_X4 U845 ( .A1(n2145), .A2(n3027), .ZN(n3125) );
  NAND2_X2 U846 ( .A1(n1764), .A2(n2092), .ZN(n1828) );
  NAND2_X2 U847 ( .A1(n3441), .A2(n1829), .ZN(n1764) );
  OAI21_X2 U848 ( .B1(n3204), .B2(n213), .A(n17), .ZN(n497) );
  INV_X2 U849 ( .A(a[3]), .ZN(n213) );
  INV_X4 U850 ( .A(n3025), .ZN(n1069) );
  NAND2_X2 U852 ( .A1(n3093), .A2(n1222), .ZN(n1428) );
  AOI22_X2 U853 ( .A1(n2228), .A2(n3200), .B1(n93), .B2(n3453), .ZN(n861) );
  INV_X4 U854 ( .A(n2111), .ZN(n1856) );
  NAND2_X4 U855 ( .A1(n1399), .A2(n1398), .ZN(n3050) );
  NAND2_X2 U856 ( .A1(n215), .A2(n214), .ZN(n1609) );
  INV_X2 U857 ( .A(n1759), .ZN(n214) );
  INV_X2 U858 ( .A(n240), .ZN(n215) );
  INV_X2 U859 ( .A(n2944), .ZN(n217) );
  NOR2_X2 U860 ( .A1(n2911), .A2(n2910), .ZN(n2944) );
  NAND3_X2 U861 ( .A1(n1482), .A2(n3999), .A3(n1892), .ZN(n3991) );
  NAND2_X2 U862 ( .A1(n3299), .A2(n3966), .ZN(n434) );
  NOR2_X2 U865 ( .A1(n1141), .A2(n1857), .ZN(n219) );
  NAND2_X2 U867 ( .A1(n2651), .A2(n1267), .ZN(n1269) );
  NAND2_X2 U868 ( .A1(n1377), .A2(n2407), .ZN(n2449) );
  NAND3_X1 U869 ( .A1(n2519), .A2(n2520), .A3(n725), .ZN(n1558) );
  NOR2_X2 U870 ( .A1(n221), .A2(n1691), .ZN(n1924) );
  INV_X4 U872 ( .A(n2327), .ZN(n2009) );
  NAND2_X2 U873 ( .A1(n2527), .A2(n1541), .ZN(n1355) );
  NOR2_X2 U874 ( .A1(n2018), .A2(n2559), .ZN(n1991) );
  INV_X4 U875 ( .A(n2741), .ZN(n585) );
  NAND3_X2 U876 ( .A1(n2677), .A2(n2676), .A3(n2678), .ZN(n809) );
  NOR2_X2 U877 ( .A1(n3204), .A2(n3413), .ZN(n2833) );
  NAND2_X2 U878 ( .A1(n3329), .A2(n37), .ZN(n2537) );
  NAND3_X2 U879 ( .A1(n896), .A2(n2575), .A3(n895), .ZN(n2631) );
  NAND2_X2 U880 ( .A1(n926), .A2(n925), .ZN(n1383) );
  NAND2_X2 U882 ( .A1(n2007), .A2(n3564), .ZN(n3565) );
  NAND2_X2 U883 ( .A1(n1715), .A2(n4056), .ZN(n2551) );
  NOR2_X2 U886 ( .A1(n76), .A2(n2285), .ZN(n2986) );
  OAI21_X2 U888 ( .B1(n3258), .B2(n3257), .A(n3281), .ZN(n385) );
  NAND2_X2 U889 ( .A1(n3255), .A2(n540), .ZN(n386) );
  NAND2_X2 U890 ( .A1(n3235), .A2(n3234), .ZN(n3236) );
  NAND2_X2 U891 ( .A1(n650), .A2(n1882), .ZN(n3235) );
  NAND2_X2 U892 ( .A1(n1474), .A2(n3021), .ZN(n1935) );
  NAND2_X2 U893 ( .A1(n224), .A2(n1573), .ZN(\d[31]_BAR ) );
  NAND2_X2 U894 ( .A1(n1571), .A2(n1572), .ZN(n224) );
  INV_X4 U895 ( .A(n2890), .ZN(n317) );
  INV_X4 U896 ( .A(n225), .ZN(n1614) );
  NOR2_X2 U897 ( .A1(n3225), .A2(n2126), .ZN(n225) );
  INV_X4 U898 ( .A(n3268), .ZN(n1900) );
  AOI21_X2 U899 ( .B1(n2385), .B2(n1265), .A(n3046), .ZN(n1831) );
  AOI21_X2 U900 ( .B1(n1486), .B2(n415), .A(n1069), .ZN(n3046) );
  INV_X4 U901 ( .A(n688), .ZN(n2544) );
  NAND3_X2 U903 ( .A1(n4018), .A2(n4019), .A3(n4017), .ZN(n4022) );
  NAND2_X2 U904 ( .A1(n1418), .A2(n2117), .ZN(n1590) );
  NAND2_X2 U905 ( .A1(n1121), .A2(a[12]), .ZN(n914) );
  INV_X8 U906 ( .A(n3009), .ZN(n249) );
  NOR2_X2 U907 ( .A1(n3204), .A2(n3016), .ZN(n2065) );
  NOR2_X2 U908 ( .A1(n3329), .A2(n205), .ZN(n2153) );
  NAND2_X2 U909 ( .A1(n226), .A2(n3172), .ZN(n975) );
  NAND2_X2 U910 ( .A1(n3170), .A2(n3171), .ZN(n226) );
  NOR2_X2 U911 ( .A1(n3177), .A2(a[7]), .ZN(n2778) );
  NOR2_X4 U912 ( .A1(b[11]), .A2(b[12]), .ZN(n1087) );
  OAI21_X2 U913 ( .B1(n3800), .B2(n3819), .A(n1312), .ZN(n3802) );
  NAND2_X2 U914 ( .A1(n1590), .A2(n1502), .ZN(n3747) );
  AOI22_X2 U915 ( .A1(n248), .A2(n2778), .B1(n3409), .B2(n247), .ZN(n246) );
  OAI21_X2 U918 ( .B1(n3558), .B2(n3805), .A(n866), .ZN(n2196) );
  NAND2_X2 U919 ( .A1(n4027), .A2(n4026), .ZN(n1573) );
  NAND2_X2 U922 ( .A1(n227), .A2(n1538), .ZN(n2051) );
  INV_X8 U923 ( .A(n1449), .ZN(n831) );
  AOI21_X2 U924 ( .B1(n2299), .B2(a[11]), .A(n3176), .ZN(n1100) );
  NAND3_X2 U927 ( .A1(n3461), .A2(n1660), .A3(n228), .ZN(n3467) );
  INV_X1 U928 ( .A(n1370), .ZN(n230) );
  INV_X2 U929 ( .A(n3734), .ZN(n1363) );
  INV_X4 U930 ( .A(n2198), .ZN(n1337) );
  NAND2_X2 U932 ( .A1(n233), .A2(n232), .ZN(n231) );
  INV_X2 U933 ( .A(n872), .ZN(n232) );
  NOR2_X2 U935 ( .A1(n4174), .A2(n4076), .ZN(n3909) );
  NOR2_X2 U936 ( .A1(n3308), .A2(n3309), .ZN(n3334) );
  OAI21_X2 U940 ( .B1(n1897), .B2(n1896), .A(n234), .ZN(n3872) );
  AOI22_X2 U941 ( .A1(n1894), .A2(n1895), .B1(n1309), .B2(n3710), .ZN(n234) );
  NAND2_X2 U942 ( .A1(n236), .A2(n235), .ZN(n2030) );
  INV_X2 U943 ( .A(n2081), .ZN(n235) );
  INV_X2 U944 ( .A(n3158), .ZN(n236) );
  XNOR2_X2 U947 ( .A(n2356), .B(n2301), .ZN(n3307) );
  NAND2_X2 U948 ( .A1(n2620), .A2(n2588), .ZN(n2587) );
  NOR2_X2 U949 ( .A1(n1337), .A2(n677), .ZN(n3137) );
  NAND3_X2 U950 ( .A1(n3712), .A2(n2061), .A3(n4021), .ZN(n3713) );
  NOR2_X4 U951 ( .A1(n641), .A2(n1983), .ZN(n4021) );
  NAND2_X2 U953 ( .A1(n1420), .A2(n1419), .ZN(n1881) );
  AOI21_X2 U954 ( .B1(n76), .B2(n2285), .A(n2994), .ZN(n2987) );
  NAND2_X2 U955 ( .A1(n4011), .A2(n1618), .ZN(n237) );
  NAND2_X2 U956 ( .A1(n662), .A2(n3133), .ZN(n1785) );
  NAND2_X2 U957 ( .A1(n1852), .A2(n1223), .ZN(n662) );
  NAND2_X2 U958 ( .A1(n1769), .A2(n3388), .ZN(n3398) );
  INV_X8 U959 ( .A(n2335), .ZN(n3454) );
  NAND3_X2 U960 ( .A1(n2336), .A2(b[4]), .A3(n2785), .ZN(n2335) );
  INV_X4 U961 ( .A(n922), .ZN(n1407) );
  NAND2_X2 U962 ( .A1(n3472), .A2(n56), .ZN(n859) );
  NAND2_X2 U963 ( .A1(n2356), .A2(n2022), .ZN(n2981) );
  NAND3_X2 U966 ( .A1(n3636), .A2(n4021), .A3(n3864), .ZN(n239) );
  NAND3_X2 U968 ( .A1(n1910), .A2(n1911), .A3(n401), .ZN(n1909) );
  NOR2_X2 U969 ( .A1(n411), .A2(n3283), .ZN(n3289) );
  NAND2_X2 U970 ( .A1(n1386), .A2(n1385), .ZN(n411) );
  NOR2_X2 U972 ( .A1(n249), .A2(n1837), .ZN(n248) );
  NOR2_X2 U973 ( .A1(n2924), .A2(n2165), .ZN(n247) );
  AOI22_X2 U974 ( .A1(n3010), .A2(n2870), .B1(n2871), .B2(n2924), .ZN(n2890)
         );
  NAND2_X1 U975 ( .A1(n240), .A2(n1759), .ZN(n1608) );
  NAND2_X2 U976 ( .A1(n306), .A2(n305), .ZN(n240) );
  MUX2_X2 U979 ( .A(n241), .B(n117), .S(a[17]), .Z(n2577) );
  MUX2_X2 U980 ( .A(n105), .B(n117), .S(a[20]), .Z(n2719) );
  MUX2_X2 U981 ( .A(n105), .B(n117), .S(n97), .Z(n2638) );
  MUX2_X2 U982 ( .A(n105), .B(n1834), .S(a[22]), .Z(n2682) );
  NAND2_X2 U983 ( .A1(n242), .A2(n499), .ZN(n3753) );
  NAND2_X2 U984 ( .A1(n1607), .A2(n1606), .ZN(n242) );
  NAND2_X2 U985 ( .A1(n726), .A2(n502), .ZN(n1606) );
  AOI22_X2 U986 ( .A1(n1661), .A2(n2263), .B1(n509), .B2(n1711), .ZN(n502) );
  BUF_X4 U989 ( .A(n2857), .Z(n244) );
  OAI21_X2 U990 ( .B1(n92), .B2(n2779), .A(n246), .ZN(n2925) );
  INV_X2 U991 ( .A(n250), .ZN(n554) );
  NAND2_X2 U992 ( .A1(n2305), .A2(n3248), .ZN(n250) );
  AOI21_X2 U993 ( .B1(n250), .B2(n768), .A(n1132), .ZN(n2146) );
  INV_X2 U996 ( .A(n253), .ZN(n252) );
  NAND2_X2 U997 ( .A1(n3792), .A2(n3561), .ZN(n3746) );
  NOR2_X2 U998 ( .A1(n2166), .A2(n3096), .ZN(n3792) );
  INV_X2 U1000 ( .A(n1627), .ZN(n546) );
  NAND2_X1 U1001 ( .A1(n3240), .A2(n1630), .ZN(n254) );
  NOR2_X2 U1002 ( .A1(n3239), .A2(n3238), .ZN(n3240) );
  NAND3_X2 U1004 ( .A1(n1952), .A2(n1948), .A3(n1949), .ZN(n1208) );
  AOI22_X2 U1005 ( .A1(n2359), .A2(n2438), .B1(n524), .B2(a[14]), .ZN(n2851)
         );
  NAND2_X2 U1007 ( .A1(n256), .A2(n255), .ZN(n793) );
  INV_X2 U1008 ( .A(n2851), .ZN(n255) );
  NAND3_X2 U1009 ( .A1(n1920), .A2(n2849), .A3(n504), .ZN(n257) );
  NAND2_X2 U1011 ( .A1(n1920), .A2(n2849), .ZN(n2850) );
  NAND3_X2 U1012 ( .A1(n258), .A2(n1632), .A3(n1789), .ZN(n4004) );
  INV_X2 U1015 ( .A(n2280), .ZN(n259) );
  NAND2_X2 U1016 ( .A1(n771), .A2(n3296), .ZN(n2280) );
  NOR2_X2 U1018 ( .A1(n2507), .A2(n264), .ZN(n261) );
  NAND2_X2 U1020 ( .A1(n4042), .A2(n2257), .ZN(n264) );
  INV_X2 U1021 ( .A(n687), .ZN(n2545) );
  INV_X2 U1022 ( .A(n265), .ZN(n266) );
  INV_X2 U1024 ( .A(n3515), .ZN(n1752) );
  XNOR2_X2 U1025 ( .A(n2907), .B(n2924), .ZN(n267) );
  AOI22_X2 U1026 ( .A1(n1360), .A2(n268), .B1(n1227), .B2(n15), .ZN(n2112) );
  INV_X2 U1027 ( .A(n269), .ZN(n268) );
  AOI22_X2 U1028 ( .A1(n2982), .A2(n2438), .B1(n3202), .B2(n3176), .ZN(n269)
         );
  INV_X4 U1029 ( .A(n1227), .ZN(n1360) );
  NOR2_X4 U1030 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  NOR2_X2 U1031 ( .A1(n272), .A2(n271), .ZN(n3253) );
  INV_X4 U1032 ( .A(n270), .ZN(n3254) );
  NAND2_X2 U1033 ( .A1(n271), .A2(n272), .ZN(n270) );
  NAND2_X2 U1034 ( .A1(n2554), .A2(n2553), .ZN(n271) );
  NAND2_X2 U1036 ( .A1(n2945), .A2(n276), .ZN(n273) );
  INV_X2 U1037 ( .A(n275), .ZN(n274) );
  INV_X2 U1038 ( .A(n1630), .ZN(n3276) );
  NAND2_X2 U1039 ( .A1(n1518), .A2(n1629), .ZN(n1630) );
  OAI22_X2 U1041 ( .A1(n278), .A2(n92), .B1(n277), .B2(n2997), .ZN(n1362) );
  AOI22_X2 U1042 ( .A1(n3139), .A2(n3034), .B1(n3177), .B2(n3413), .ZN(n277)
         );
  INV_X2 U1043 ( .A(n2521), .ZN(n1307) );
  NAND2_X2 U1044 ( .A1(n2519), .A2(n2520), .ZN(n2521) );
  NAND2_X1 U1045 ( .A1(n2440), .A2(n1898), .ZN(n2520) );
  NAND2_X2 U1047 ( .A1(n280), .A2(n279), .ZN(n2519) );
  NAND2_X2 U1049 ( .A1(n281), .A2(n2066), .ZN(n1570) );
  NAND2_X2 U1050 ( .A1(n281), .A2(n1311), .ZN(n3979) );
  NAND3_X2 U1051 ( .A1(n2066), .A2(n3710), .A3(n281), .ZN(n1897) );
  NAND2_X2 U1052 ( .A1(n60), .A2(n1409), .ZN(n281) );
  INV_X1 U1055 ( .A(n3959), .ZN(n284) );
  INV_X1 U1056 ( .A(n1991), .ZN(n2525) );
  INV_X2 U1057 ( .A(n724), .ZN(n723) );
  NAND2_X2 U1058 ( .A1(n289), .A2(n285), .ZN(n724) );
  NAND2_X2 U1059 ( .A1(n288), .A2(n286), .ZN(n285) );
  NOR2_X2 U1060 ( .A1(n287), .A2(n1991), .ZN(n286) );
  INV_X1 U1061 ( .A(n2524), .ZN(n287) );
  NAND2_X2 U1062 ( .A1(n2547), .A2(n2530), .ZN(n288) );
  NAND2_X2 U1063 ( .A1(n290), .A2(n2529), .ZN(n289) );
  NAND3_X2 U1064 ( .A1(n2531), .A2(n2530), .A3(n1991), .ZN(n290) );
  INV_X4 U1065 ( .A(n2785), .ZN(n2145) );
  NAND2_X2 U1066 ( .A1(n1024), .A2(n1023), .ZN(n857) );
  NAND2_X1 U1067 ( .A1(b[6]), .A2(n2334), .ZN(n1023) );
  INV_X2 U1068 ( .A(b[6]), .ZN(n291) );
  NAND2_X2 U1069 ( .A1(n292), .A2(n4161), .ZN(n1445) );
  INV_X2 U1070 ( .A(n2368), .ZN(n292) );
  NAND3_X2 U1071 ( .A1(n1772), .A2(n3706), .A3(n3705), .ZN(\d[32] ) );
  OAI22_X2 U1072 ( .A1(n3835), .A2(n3834), .B1(n293), .B2(n3836), .ZN(\d[18] )
         );
  NOR2_X2 U1074 ( .A1(n297), .A2(n295), .ZN(n3905) );
  NAND2_X2 U1075 ( .A1(n294), .A2(n3820), .ZN(n3828) );
  INV_X2 U1076 ( .A(n297), .ZN(n294) );
  NAND2_X2 U1077 ( .A1(n296), .A2(n3820), .ZN(n295) );
  NOR2_X2 U1079 ( .A1(n2090), .A2(n3791), .ZN(n297) );
  NOR2_X2 U1081 ( .A1(n3313), .A2(n3312), .ZN(n3385) );
  NAND2_X2 U1083 ( .A1(n831), .A2(n99), .ZN(n300) );
  NAND2_X2 U1084 ( .A1(n302), .A2(n3704), .ZN(n3706) );
  NAND2_X2 U1085 ( .A1(n3695), .A2(n302), .ZN(n3696) );
  NAND2_X2 U1086 ( .A1(n3631), .A2(n302), .ZN(n3634) );
  NOR3_X2 U1087 ( .A1(n302), .A2(n3635), .A3(n181), .ZN(n3624) );
  NOR2_X4 U1088 ( .A1(n1288), .A2(n1363), .ZN(n302) );
  NAND2_X2 U1089 ( .A1(n304), .A2(n303), .ZN(n1759) );
  NAND2_X2 U1091 ( .A1(n65), .A2(n334), .ZN(n304) );
  NAND2_X2 U1092 ( .A1(n1758), .A2(n3086), .ZN(n306) );
  NOR2_X2 U1094 ( .A1(n902), .A2(n307), .ZN(n901) );
  NAND2_X2 U1095 ( .A1(n1702), .A2(n307), .ZN(n898) );
  INV_X4 U1096 ( .A(n312), .ZN(n307) );
  NAND2_X2 U1097 ( .A1(n309), .A2(n308), .ZN(n1504) );
  INV_X2 U1098 ( .A(n2965), .ZN(n308) );
  AOI21_X2 U1099 ( .B1(n2928), .B2(n2929), .A(n2927), .ZN(n2965) );
  NOR2_X2 U1100 ( .A1(n2839), .A2(n2840), .ZN(n2927) );
  NAND2_X2 U1101 ( .A1(n2840), .A2(n2839), .ZN(n2929) );
  NOR2_X2 U1102 ( .A1(n2843), .A2(n2842), .ZN(n2928) );
  NAND2_X2 U1103 ( .A1(n1076), .A2(n1959), .ZN(n309) );
  NAND2_X2 U1105 ( .A1(n311), .A2(n310), .ZN(n1076) );
  INV_X2 U1106 ( .A(n2963), .ZN(n310) );
  NAND2_X2 U1108 ( .A1(n2140), .A2(n2141), .ZN(n311) );
  NAND2_X2 U1109 ( .A1(n2142), .A2(n2953), .ZN(n2141) );
  NAND3_X2 U1111 ( .A1(n2977), .A2(n312), .A3(n1702), .ZN(n1701) );
  NAND2_X2 U1113 ( .A1(n2161), .A2(n426), .ZN(n315) );
  NAND2_X2 U1114 ( .A1(n318), .A2(n317), .ZN(n316) );
  INV_X2 U1115 ( .A(n2271), .ZN(n319) );
  BUF_X4 U1116 ( .A(n3034), .Z(n313) );
  NAND2_X2 U1117 ( .A1(n2880), .A2(n314), .ZN(n1832) );
  NAND2_X2 U1118 ( .A1(n316), .A2(n315), .ZN(n2880) );
  NAND2_X2 U1119 ( .A1(n319), .A2(n3034), .ZN(n318) );
  INV_X2 U1124 ( .A(n2564), .ZN(n2562) );
  INV_X2 U1125 ( .A(n324), .ZN(n2563) );
  INV_X4 U1127 ( .A(n1448), .ZN(n3120) );
  INV_X4 U1128 ( .A(n1302), .ZN(n3119) );
  INV_X2 U1129 ( .A(n2420), .ZN(n2417) );
  NAND2_X2 U1130 ( .A1(n328), .A2(n325), .ZN(n2420) );
  NOR2_X1 U1131 ( .A1(n2411), .A2(n3128), .ZN(n326) );
  INV_X2 U1133 ( .A(n329), .ZN(n328) );
  NOR2_X2 U1134 ( .A1(n2413), .A2(n330), .ZN(n329) );
  XNOR2_X2 U1135 ( .A(n2740), .B(n3124), .ZN(n330) );
  NOR2_X2 U1136 ( .A1(n384), .A2(n1510), .ZN(n3299) );
  NOR2_X4 U1137 ( .A1(n674), .A2(n1395), .ZN(n1510) );
  NAND2_X2 U1138 ( .A1(n3978), .A2(n4003), .ZN(n384) );
  BUF_X4 U1139 ( .A(n3087), .Z(n333) );
  INV_X2 U1140 ( .A(n3087), .ZN(n334) );
  INV_X2 U1143 ( .A(n1492), .ZN(n336) );
  OAI21_X2 U1144 ( .B1(n338), .B2(n1492), .A(n3380), .ZN(n337) );
  INV_X2 U1145 ( .A(n3381), .ZN(n338) );
  NAND2_X2 U1146 ( .A1(n839), .A2(n2671), .ZN(n3381) );
  NAND2_X2 U1147 ( .A1(n339), .A2(a[13]), .ZN(n2849) );
  NAND2_X2 U1148 ( .A1(n339), .A2(a[17]), .ZN(n1930) );
  AOI22_X1 U1149 ( .A1(n1863), .A2(n2697), .B1(n339), .B2(a[22]), .ZN(n356) );
  INV_X2 U1150 ( .A(n4075), .ZN(n339) );
  NAND2_X2 U1153 ( .A1(n1932), .A2(n402), .ZN(n340) );
  NAND2_X2 U1154 ( .A1(n343), .A2(n341), .ZN(n1265) );
  NAND3_X2 U1155 ( .A1(n342), .A2(n1932), .A3(n402), .ZN(n341) );
  INV_X2 U1156 ( .A(n344), .ZN(n342) );
  INV_X1 U1157 ( .A(n3183), .ZN(n969) );
  AOI21_X2 U1158 ( .B1(n608), .B2(n3199), .A(n607), .ZN(n401) );
  NOR2_X2 U1159 ( .A1(n1223), .A2(n347), .ZN(n607) );
  XNOR2_X2 U1160 ( .A(n345), .B(n346), .ZN(n3199) );
  XNOR2_X2 U1161 ( .A(n1116), .B(n3183), .ZN(n345) );
  NAND3_X2 U1162 ( .A1(n796), .A2(n1117), .A3(n795), .ZN(n1116) );
  NOR2_X2 U1163 ( .A1(n3181), .A2(n3182), .ZN(n346) );
  INV_X2 U1165 ( .A(n3198), .ZN(n347) );
  AOI21_X2 U1166 ( .B1(n4065), .B2(n1046), .A(n3135), .ZN(n3198) );
  NAND2_X2 U1167 ( .A1(n3220), .A2(n412), .ZN(n1342) );
  OAI21_X2 U1170 ( .B1(n1875), .B2(n2106), .A(n1286), .ZN(n837) );
  NAND2_X2 U1171 ( .A1(n1855), .A2(n2721), .ZN(n838) );
  NAND2_X2 U1174 ( .A1(n75), .A2(n842), .ZN(n349) );
  NAND3_X1 U1175 ( .A1(n1014), .A2(n350), .A3(n1013), .ZN(n1275) );
  NAND2_X2 U1176 ( .A1(n1683), .A2(n2973), .ZN(n1013) );
  INV_X2 U1177 ( .A(n2974), .ZN(n350) );
  NAND2_X2 U1179 ( .A1(n1680), .A2(n2858), .ZN(n351) );
  NAND2_X2 U1180 ( .A1(n574), .A2(n2860), .ZN(n352) );
  NAND2_X2 U1181 ( .A1(n72), .A2(n1595), .ZN(n1014) );
  INV_X4 U1182 ( .A(n1683), .ZN(n1595) );
  NAND2_X4 U1184 ( .A1(n1682), .A2(n1681), .ZN(n2973) );
  NAND3_X2 U1185 ( .A1(n355), .A2(n354), .A3(n353), .ZN(n2110) );
  NAND2_X2 U1186 ( .A1(n2737), .A2(n3109), .ZN(n353) );
  NAND2_X2 U1188 ( .A1(n357), .A2(n356), .ZN(n688) );
  NAND2_X2 U1189 ( .A1(n1645), .A2(n445), .ZN(n357) );
  BUF_X4 U1190 ( .A(n1102), .Z(n358) );
  NOR2_X2 U1195 ( .A1(n1697), .A2(n3290), .ZN(n360) );
  INV_X2 U1197 ( .A(n424), .ZN(n362) );
  NAND2_X2 U1198 ( .A1(n376), .A2(n2128), .ZN(n363) );
  NAND2_X2 U1199 ( .A1(n365), .A2(n364), .ZN(n2147) );
  NAND2_X1 U1200 ( .A1(n2146), .A2(n3297), .ZN(n364) );
  XNOR2_X2 U1202 ( .A(n1440), .B(n366), .ZN(n3284) );
  NAND2_X2 U1204 ( .A1(n3291), .A2(n1102), .ZN(n370) );
  NAND2_X2 U1206 ( .A1(n2544), .A2(n2545), .ZN(n372) );
  NOR2_X2 U1207 ( .A1(n1367), .A2(n447), .ZN(n371) );
  NAND2_X2 U1208 ( .A1(n687), .A2(n688), .ZN(n373) );
  INV_X4 U1209 ( .A(n374), .ZN(n1989) );
  NAND2_X2 U1210 ( .A1(n1902), .A2(n1899), .ZN(n374) );
  NAND2_X2 U1214 ( .A1(n1988), .A2(n1987), .ZN(n375) );
  INV_X2 U1215 ( .A(n3284), .ZN(n1985) );
  INV_X2 U1216 ( .A(n3285), .ZN(n1986) );
  NAND2_X2 U1217 ( .A1(n1989), .A2(n1984), .ZN(n3956) );
  NAND2_X2 U1218 ( .A1(n3285), .A2(n3284), .ZN(n1987) );
  INV_X4 U1220 ( .A(n1697), .ZN(n376) );
  NAND2_X2 U1222 ( .A1(n2127), .A2(n378), .ZN(n382) );
  INV_X4 U1223 ( .A(n3270), .ZN(n378) );
  NOR2_X2 U1224 ( .A1(n719), .A2(n718), .ZN(n717) );
  NAND2_X2 U1225 ( .A1(n380), .A2(n379), .ZN(n718) );
  NAND2_X2 U1226 ( .A1(n1939), .A2(n3288), .ZN(n379) );
  NAND2_X2 U1227 ( .A1(n383), .A2(n1440), .ZN(n380) );
  INV_X2 U1229 ( .A(n1697), .ZN(n1539) );
  NOR2_X2 U1230 ( .A1(n3270), .A2(n3269), .ZN(n3286) );
  NAND2_X2 U1231 ( .A1(n377), .A2(n376), .ZN(n381) );
  NAND2_X2 U1232 ( .A1(n3273), .A2(n3272), .ZN(n3288) );
  INV_X2 U1233 ( .A(n1939), .ZN(n383) );
  NAND2_X2 U1236 ( .A1(n1366), .A2(n1367), .ZN(n388) );
  INV_X2 U1237 ( .A(n2528), .ZN(n744) );
  INV_X4 U1238 ( .A(n1870), .ZN(n2500) );
  NAND2_X2 U1239 ( .A1(n391), .A2(n390), .ZN(n2447) );
  OAI22_X2 U1240 ( .A1(n2246), .A2(n2245), .B1(n2488), .B2(n2486), .ZN(n390)
         );
  AOI21_X2 U1241 ( .B1(n393), .B2(n2446), .A(n392), .ZN(n2448) );
  NOR2_X2 U1242 ( .A1(n1686), .A2(n742), .ZN(n392) );
  NAND2_X1 U1243 ( .A1(n742), .A2(n1686), .ZN(n393) );
  INV_X2 U1244 ( .A(n3267), .ZN(n1903) );
  NAND2_X2 U1245 ( .A1(n936), .A2(n935), .ZN(n3267) );
  NAND2_X2 U1246 ( .A1(n395), .A2(n394), .ZN(n935) );
  NAND2_X2 U1247 ( .A1(n2160), .A2(n2568), .ZN(n394) );
  NAND2_X2 U1248 ( .A1(n1403), .A2(n1404), .ZN(n395) );
  NAND2_X2 U1249 ( .A1(n397), .A2(n396), .ZN(n936) );
  NAND3_X2 U1250 ( .A1(n1169), .A2(n2208), .A3(n2207), .ZN(n396) );
  NAND2_X2 U1251 ( .A1(n2159), .A2(n1354), .ZN(n397) );
  INV_X2 U1252 ( .A(n1866), .ZN(n1865) );
  INV_X2 U1253 ( .A(n1869), .ZN(n1868) );
  NAND2_X2 U1254 ( .A1(n399), .A2(n1867), .ZN(n1329) );
  NAND3_X2 U1255 ( .A1(n2115), .A2(n1123), .A3(n2114), .ZN(n1867) );
  NOR2_X2 U1256 ( .A1(n1869), .A2(n1866), .ZN(n399) );
  NOR2_X2 U1258 ( .A1(n1911), .A2(n401), .ZN(n609) );
  NAND2_X4 U1260 ( .A1(n1645), .A2(n440), .ZN(n402) );
  NAND2_X2 U1264 ( .A1(n2844), .A2(n2928), .ZN(n403) );
  NAND2_X2 U1265 ( .A1(n1476), .A2(n1477), .ZN(n404) );
  NAND2_X4 U1266 ( .A1(n406), .A2(n405), .ZN(n1300) );
  NAND2_X2 U1271 ( .A1(n1904), .A2(n409), .ZN(n722) );
  OAI21_X2 U1272 ( .B1(n1557), .B2(n4141), .A(n73), .ZN(n409) );
  NAND2_X2 U1273 ( .A1(n410), .A2(n2974), .ZN(n1274) );
  NAND2_X2 U1274 ( .A1(n1014), .A2(n1013), .ZN(n410) );
  NAND2_X2 U1276 ( .A1(n3222), .A2(n3221), .ZN(n412) );
  INV_X2 U1277 ( .A(n415), .ZN(n490) );
  OAI21_X2 U1278 ( .B1(n1069), .B2(n1070), .A(n415), .ZN(n870) );
  NAND2_X2 U1284 ( .A1(n418), .A2(n3382), .ZN(n3803) );
  NAND2_X2 U1285 ( .A1(n3338), .A2(n3337), .ZN(n3382) );
  NAND2_X2 U1286 ( .A1(n419), .A2(n3383), .ZN(n418) );
  NAND2_X2 U1287 ( .A1(n3335), .A2(n3336), .ZN(n3383) );
  NAND4_X1 U1288 ( .A1(n823), .A2(n821), .A3(n4140), .A4(n824), .ZN(n419) );
  NAND3_X2 U1289 ( .A1(n422), .A2(n49), .A3(n420), .ZN(n714) );
  NAND2_X1 U1290 ( .A1(n1659), .A2(a[8]), .ZN(n420) );
  NAND2_X2 U1295 ( .A1(n1375), .A2(n1376), .ZN(n425) );
  NAND2_X2 U1296 ( .A1(n1375), .A2(n1376), .ZN(n930) );
  INV_X4 U1297 ( .A(n2919), .ZN(n773) );
  NAND2_X4 U1298 ( .A1(n503), .A2(n2229), .ZN(n3058) );
  INV_X4 U1299 ( .A(n1786), .ZN(n644) );
  INV_X1 U1300 ( .A(n2880), .ZN(n1602) );
  INV_X1 U1302 ( .A(n3725), .ZN(n3712) );
  NAND2_X2 U1303 ( .A1(n1498), .A2(n3103), .ZN(n1364) );
  NAND2_X4 U1304 ( .A1(n1038), .A2(n3171), .ZN(n3228) );
  NOR2_X1 U1306 ( .A1(n4051), .A2(n2193), .ZN(n749) );
  NAND2_X2 U1309 ( .A1(n938), .A2(n937), .ZN(n2529) );
  OAI21_X1 U1312 ( .B1(n1298), .B2(n3050), .A(n3049), .ZN(n431) );
  NAND2_X2 U1313 ( .A1(n1024), .A2(n1023), .ZN(n432) );
  NAND2_X4 U1314 ( .A1(n2009), .A2(n2326), .ZN(n2329) );
  INV_X4 U1318 ( .A(n1301), .ZN(n1302) );
  NAND2_X4 U1319 ( .A1(n3990), .A2(n2247), .ZN(n951) );
  INV_X1 U1320 ( .A(n925), .ZN(n594) );
  NAND2_X1 U1321 ( .A1(n3948), .A2(n3949), .ZN(n3952) );
  NAND2_X1 U1322 ( .A1(n1455), .A2(n1456), .ZN(n1458) );
  NAND2_X1 U1323 ( .A1(n1456), .A2(n2985), .ZN(n1703) );
  NOR2_X2 U1324 ( .A1(n2983), .A2(n463), .ZN(n3136) );
  NOR2_X4 U1325 ( .A1(n1780), .A2(n1783), .ZN(n2018) );
  NOR3_X4 U1327 ( .A1(n1323), .A2(b[8]), .A3(b[7]), .ZN(n1845) );
  NAND2_X1 U1328 ( .A1(n3225), .A2(n2126), .ZN(n1613) );
  NOR2_X2 U1329 ( .A1(n3303), .A2(a[10]), .ZN(n1099) );
  NOR2_X4 U1330 ( .A1(n1727), .A2(n1726), .ZN(n3059) );
  NAND2_X2 U1331 ( .A1(n1397), .A2(n3467), .ZN(n1278) );
  NOR3_X1 U1333 ( .A1(n3940), .A2(n3936), .A3(n4005), .ZN(n3935) );
  NOR2_X2 U1334 ( .A1(n3605), .A2(n1363), .ZN(n3863) );
  NAND2_X2 U1335 ( .A1(n617), .A2(n2018), .ZN(n1443) );
  NOR2_X1 U1336 ( .A1(n2850), .A2(n2851), .ZN(n673) );
  NAND2_X2 U1337 ( .A1(n425), .A2(n929), .ZN(n437) );
  NAND3_X1 U1339 ( .A1(n2412), .A2(n2316), .A3(n1315), .ZN(n2411) );
  NAND2_X1 U1340 ( .A1(n3981), .A2(n2286), .ZN(n3895) );
  OAI21_X2 U1341 ( .B1(n804), .B2(n803), .A(n802), .ZN(n1635) );
  INV_X4 U1342 ( .A(n2829), .ZN(n803) );
  INV_X1 U1343 ( .A(n2977), .ZN(n902) );
  NOR2_X4 U1344 ( .A1(n2930), .A2(n2931), .ZN(n2138) );
  NAND2_X2 U1345 ( .A1(n3241), .A2(n2063), .ZN(n1625) );
  INV_X2 U1346 ( .A(n2138), .ZN(n1349) );
  NOR2_X2 U1347 ( .A1(n87), .A2(a[20]), .ZN(n2549) );
  AOI22_X2 U1348 ( .A1(n3034), .A2(a[7]), .B1(n249), .B2(n3468), .ZN(n2779) );
  NOR2_X1 U1349 ( .A1(n3642), .A2(n3840), .ZN(n3844) );
  NOR2_X1 U1350 ( .A1(n3123), .A2(n2441), .ZN(n1120) );
  NAND2_X2 U1351 ( .A1(n3113), .A2(a[8]), .ZN(n1854) );
  NAND2_X2 U1352 ( .A1(n3839), .A2(n3413), .ZN(n3114) );
  NOR2_X1 U1353 ( .A1(n2907), .A2(a[12]), .ZN(n2414) );
  NOR2_X1 U1354 ( .A1(n3016), .A2(b[14]), .ZN(n2415) );
  NAND2_X1 U1355 ( .A1(n1362), .A2(n3149), .ZN(n3150) );
  INV_X1 U1356 ( .A(n2957), .ZN(n2958) );
  NOR2_X2 U1358 ( .A1(n3144), .A2(n3180), .ZN(n3158) );
  NAND2_X1 U1359 ( .A1(n3055), .A2(n3057), .ZN(n1193) );
  MUX2_X1 U1361 ( .A(n3454), .B(n3455), .S(n3589), .Z(n2498) );
  MUX2_X2 U1362 ( .A(n85), .B(n1261), .S(a[8]), .Z(n2978) );
  INV_X1 U1363 ( .A(n3281), .ZN(n2328) );
  NOR2_X1 U1364 ( .A1(n79), .A2(n2635), .ZN(n2636) );
  AOI21_X1 U1365 ( .B1(n79), .B2(n2635), .A(n2634), .ZN(n2637) );
  OAI21_X1 U1367 ( .B1(n3343), .B2(n3341), .A(n3342), .ZN(n3368) );
  INV_X1 U1368 ( .A(n1021), .ZN(n3341) );
  OAI21_X1 U1369 ( .B1(n3033), .B2(n3032), .A(n4063), .ZN(n1021) );
  NAND2_X1 U1370 ( .A1(n3504), .A2(n3503), .ZN(n3509) );
  NAND2_X1 U1371 ( .A1(n1088), .A2(n2355), .ZN(n3503) );
  NAND2_X1 U1375 ( .A1(n3509), .A2(n3508), .ZN(n3521) );
  INV_X1 U1376 ( .A(n3370), .ZN(n3560) );
  NOR3_X1 U1377 ( .A1(n3654), .A2(n3653), .A3(n3652), .ZN(n3847) );
  NOR2_X1 U1378 ( .A1(n3600), .A2(n3599), .ZN(n3658) );
  INV_X2 U1381 ( .A(n4186), .ZN(n3748) );
  INV_X1 U1382 ( .A(n1823), .ZN(n1105) );
  INV_X1 U1383 ( .A(n1824), .ZN(n1106) );
  NOR2_X2 U1384 ( .A1(n2170), .A2(n2168), .ZN(n1824) );
  NOR2_X1 U1385 ( .A1(n3204), .A2(n2438), .ZN(n2168) );
  NOR2_X1 U1386 ( .A1(n1361), .A2(n55), .ZN(n2170) );
  XOR2_X1 U1387 ( .A(n3122), .B(a[15]), .Z(n2836) );
  NAND2_X1 U1388 ( .A1(n3839), .A2(n2079), .ZN(n2453) );
  AOI21_X1 U1389 ( .B1(n969), .B2(n1116), .A(n3182), .ZN(n794) );
  NAND2_X1 U1393 ( .A1(n2228), .A2(b[14]), .ZN(n2534) );
  NAND2_X1 U1394 ( .A1(n93), .A2(n2907), .ZN(n2535) );
  XNOR2_X1 U1395 ( .A(n1651), .B(a[22]), .ZN(n2425) );
  INV_X4 U1397 ( .A(n734), .ZN(n735) );
  NOR2_X1 U1398 ( .A1(n2405), .A2(n2441), .ZN(n948) );
  XNOR2_X1 U1399 ( .A(a[23]), .B(n3122), .ZN(n2405) );
  NAND2_X1 U1400 ( .A1(n4059), .A2(n1716), .ZN(n2465) );
  NAND2_X1 U1403 ( .A1(n2444), .A2(n2443), .ZN(n2445) );
  NAND2_X1 U1404 ( .A1(n3323), .A2(a[19]), .ZN(n2443) );
  XOR2_X1 U1407 ( .A(n1651), .B(a[11]), .Z(n2809) );
  NAND2_X1 U1408 ( .A1(n3177), .A2(n3139), .ZN(n3140) );
  INV_X1 U1409 ( .A(n3193), .ZN(n3196) );
  NOR2_X1 U1410 ( .A1(n3193), .A2(n1343), .ZN(n3189) );
  NAND2_X1 U1413 ( .A1(n3008), .A2(n3515), .ZN(n3011) );
  XNOR2_X1 U1415 ( .A(n3065), .B(a[12]), .ZN(n2991) );
  NAND2_X1 U1416 ( .A1(n3472), .A2(a[12]), .ZN(n2797) );
  NOR3_X2 U1419 ( .A1(n2756), .A2(n2755), .A3(n2761), .ZN(n2767) );
  AOI22_X1 U1421 ( .A1(a[20]), .A2(n1209), .B1(n1863), .B2(n3109), .ZN(n1129)
         );
  NAND2_X1 U1422 ( .A1(n1854), .A2(n3114), .ZN(n3115) );
  NOR2_X1 U1423 ( .A1(n2246), .A2(n2488), .ZN(n741) );
  INV_X1 U1424 ( .A(n2418), .ZN(n2419) );
  NAND2_X1 U1425 ( .A1(n1784), .A2(n2907), .ZN(n2823) );
  XNOR2_X1 U1426 ( .A(n3027), .B(a[12]), .ZN(n1057) );
  NAND2_X1 U1427 ( .A1(n2885), .A2(n3392), .ZN(n2886) );
  NAND2_X2 U1428 ( .A1(n2495), .A2(n2494), .ZN(n2585) );
  AOI22_X1 U1433 ( .A1(n1270), .A2(n79), .B1(n2631), .B2(n2576), .ZN(n787) );
  INV_X1 U1434 ( .A(n2576), .ZN(n1270) );
  XNOR2_X1 U1435 ( .A(n2632), .B(n2633), .ZN(n2576) );
  MUX2_X2 U1436 ( .A(n2058), .B(n155), .S(n1784), .Z(n3005) );
  NAND2_X1 U1438 ( .A1(n1121), .A2(a[11]), .ZN(n487) );
  INV_X1 U1439 ( .A(n2689), .ZN(n2690) );
  NAND3_X1 U1440 ( .A1(n1625), .A2(n1624), .A3(n3276), .ZN(n1125) );
  NAND2_X2 U1441 ( .A1(n2030), .A2(n2031), .ZN(n2036) );
  INV_X2 U1442 ( .A(n1788), .ZN(n3165) );
  XNOR2_X1 U1443 ( .A(n94), .B(n1651), .ZN(n2841) );
  NAND2_X1 U1444 ( .A1(n2915), .A2(n2916), .ZN(n670) );
  XNOR2_X1 U1445 ( .A(n3065), .B(n3124), .ZN(n2828) );
  NOR2_X1 U1446 ( .A1(n2983), .A2(n2826), .ZN(n2049) );
  NOR2_X1 U1447 ( .A1(n2907), .A2(a[1]), .ZN(n2902) );
  NOR2_X1 U1448 ( .A1(n2045), .A2(b[14]), .ZN(n2901) );
  NOR2_X1 U1449 ( .A1(n2899), .A2(n89), .ZN(n874) );
  NAND2_X1 U1450 ( .A1(n1361), .A2(n2045), .ZN(n826) );
  NAND2_X1 U1451 ( .A1(n1862), .A2(n3139), .ZN(n568) );
  XNOR2_X1 U1452 ( .A(a[1]), .B(n3498), .ZN(n3505) );
  NAND2_X1 U1453 ( .A1(n789), .A2(n787), .ZN(n2648) );
  INV_X1 U1454 ( .A(n2675), .ZN(n1433) );
  XNOR2_X1 U1455 ( .A(n2667), .B(n2668), .ZN(n2642) );
  INV_X1 U1456 ( .A(n3038), .ZN(n3041) );
  MUX2_X2 U1457 ( .A(n3455), .B(n3454), .S(n3475), .Z(n3312) );
  NAND2_X1 U1458 ( .A1(n640), .A2(n639), .ZN(n3313) );
  NAND2_X1 U1459 ( .A1(n205), .A2(n3453), .ZN(n639) );
  NAND2_X1 U1460 ( .A1(n1088), .A2(n3118), .ZN(n3035) );
  INV_X4 U1461 ( .A(n2506), .ZN(n2336) );
  NOR2_X1 U1463 ( .A1(n2441), .A2(n916), .ZN(n3532) );
  NAND2_X2 U1464 ( .A1(n3413), .A2(n1088), .ZN(n3326) );
  NAND2_X2 U1466 ( .A1(n3515), .A2(n3392), .ZN(n3394) );
  INV_X1 U1467 ( .A(n3394), .ZN(n3433) );
  NAND3_X1 U1468 ( .A1(n3370), .A2(n867), .A3(n1644), .ZN(n866) );
  OAI21_X1 U1469 ( .B1(n554), .B2(n1132), .A(n553), .ZN(n549) );
  NAND2_X2 U1470 ( .A1(n3331), .A2(n23), .ZN(n3400) );
  INV_X1 U1472 ( .A(n3889), .ZN(n890) );
  INV_X1 U1473 ( .A(n3337), .ZN(n3321) );
  NOR2_X1 U1474 ( .A1(n3597), .A2(n3596), .ZN(n3647) );
  NOR2_X1 U1475 ( .A1(n3595), .A2(n3594), .ZN(n3596) );
  AOI21_X1 U1476 ( .B1(n3595), .B2(n3594), .A(n3593), .ZN(n3597) );
  INV_X1 U1477 ( .A(n3592), .ZN(n3594) );
  NAND2_X2 U1481 ( .A1(n2289), .A2(n3746), .ZN(n2011) );
  NAND2_X1 U1482 ( .A1(n3838), .A2(n3837), .ZN(n3849) );
  MUX2_X1 U1485 ( .A(b[14]), .B(n3839), .S(n2613), .Z(n3842) );
  NOR2_X1 U1486 ( .A1(n2723), .A2(n2764), .ZN(n2724) );
  AOI21_X1 U1487 ( .B1(n2723), .B2(n2764), .A(n2768), .ZN(n2725) );
  NAND2_X1 U1488 ( .A1(n2727), .A2(n2726), .ZN(n2746) );
  OAI21_X1 U1489 ( .B1(n2730), .B2(n2729), .A(n2728), .ZN(n3580) );
  NAND2_X1 U1490 ( .A1(n3711), .A2(n14), .ZN(n3721) );
  NOR2_X1 U1491 ( .A1(n64), .A2(n10), .ZN(n751) );
  INV_X2 U1492 ( .A(n602), .ZN(n601) );
  NOR2_X1 U1494 ( .A1(n3521), .A2(n3511), .ZN(n3525) );
  INV_X1 U1495 ( .A(n3517), .ZN(n3510) );
  NAND3_X1 U1496 ( .A1(n74), .A2(n3524), .A3(n3525), .ZN(n1667) );
  NOR2_X1 U1498 ( .A1(n3798), .A2(n3809), .ZN(n3812) );
  NAND2_X1 U1500 ( .A1(n3615), .A2(n3868), .ZN(n3664) );
  NAND3_X1 U1501 ( .A1(n3967), .A2(n3987), .A3(n1617), .ZN(n3974) );
  NOR2_X1 U1502 ( .A1(n3850), .A2(n3847), .ZN(n3865) );
  NAND2_X1 U1503 ( .A1(n3664), .A2(n3663), .ZN(n3856) );
  AOI22_X1 U1504 ( .A1(n3849), .A2(n3865), .B1(n3847), .B2(n3850), .ZN(n3857)
         );
  NAND2_X1 U1505 ( .A1(n3851), .A2(n3850), .ZN(n3853) );
  INV_X1 U1506 ( .A(n3849), .ZN(n3851) );
  INV_X1 U1507 ( .A(n3721), .ZN(n3719) );
  NOR3_X2 U1509 ( .A1(n22), .A2(n3954), .A3(n3955), .ZN(n3957) );
  OR2_X1 U1513 ( .A1(n3669), .A2(n3668), .ZN(n2388) );
  NAND2_X1 U1514 ( .A1(n3813), .A2(n3812), .ZN(n3818) );
  NAND2_X1 U1515 ( .A1(n3780), .A2(n3781), .ZN(n516) );
  NOR2_X1 U1516 ( .A1(n3774), .A2(n3783), .ZN(n514) );
  NAND2_X1 U1519 ( .A1(n3752), .A2(n3754), .ZN(n3890) );
  INV_X1 U1520 ( .A(n1672), .ZN(n3768) );
  OAI21_X1 U1521 ( .B1(n3898), .B2(n3897), .A(n3896), .ZN(n3899) );
  NAND2_X1 U1522 ( .A1(n3984), .A2(n3983), .ZN(n3982) );
  AOI22_X1 U1524 ( .A1(n3997), .A2(n3999), .B1(n3998), .B2(n3996), .ZN(n4001)
         );
  NAND2_X1 U1525 ( .A1(n3830), .A2(n3826), .ZN(n3836) );
  NAND3_X1 U1526 ( .A1(n3833), .A2(n3832), .A3(n3831), .ZN(n3834) );
  NOR2_X1 U1529 ( .A1(n1621), .A2(n4005), .ZN(n4016) );
  INV_X1 U1530 ( .A(n3742), .ZN(n3740) );
  XNOR2_X1 U1531 ( .A(a[21]), .B(n1651), .ZN(n2401) );
  NAND2_X1 U1532 ( .A1(n3323), .A2(n2057), .ZN(n2536) );
  NAND2_X1 U1534 ( .A1(n96), .A2(n249), .ZN(n2075) );
  NAND2_X1 U1535 ( .A1(n3454), .A2(a[22]), .ZN(n947) );
  NAND2_X1 U1536 ( .A1(n3455), .A2(n2697), .ZN(n946) );
  NAND2_X1 U1537 ( .A1(n3472), .A2(a[23]), .ZN(n1716) );
  INV_X1 U1538 ( .A(n3146), .ZN(n3147) );
  NOR2_X1 U1539 ( .A1(n3109), .A2(n2982), .ZN(n3146) );
  OAI21_X1 U1540 ( .B1(a[20]), .B2(n2982), .A(a[21]), .ZN(n677) );
  AOI21_X1 U1542 ( .B1(n1720), .B2(n3407), .A(n448), .ZN(n979) );
  INV_X4 U1543 ( .A(n2298), .ZN(n2777) );
  NOR2_X1 U1547 ( .A1(n4075), .A2(n3217), .ZN(n1738) );
  NAND3_X1 U1548 ( .A1(n80), .A2(n1824), .A3(n1823), .ZN(n1103) );
  NAND2_X1 U1549 ( .A1(n2982), .A2(a[25]), .ZN(n2434) );
  OAI21_X1 U1550 ( .B1(n3329), .B2(a[17]), .A(n2389), .ZN(n2505) );
  NAND2_X1 U1551 ( .A1(n3839), .A2(n2258), .ZN(n2257) );
  NAND2_X1 U1553 ( .A1(n3454), .A2(n96), .ZN(n2838) );
  NAND2_X2 U1554 ( .A1(n1776), .A2(n1775), .ZN(n1045) );
  NAND2_X1 U1556 ( .A1(n3202), .A2(n2145), .ZN(n2786) );
  XOR2_X1 U1557 ( .A(n3122), .B(a[14]), .Z(n2788) );
  OAI21_X1 U1558 ( .B1(n3202), .B2(n2802), .A(n3065), .ZN(n2217) );
  AOI22_X1 U1559 ( .A1(n3176), .A2(n3128), .B1(n2400), .B2(n2982), .ZN(n2872)
         );
  NOR2_X1 U1560 ( .A1(n2028), .A2(n3010), .ZN(n2027) );
  NOR2_X1 U1561 ( .A1(n1890), .A2(n55), .ZN(n1889) );
  NAND2_X1 U1562 ( .A1(n1818), .A2(n3128), .ZN(n3130) );
  NAND2_X1 U1563 ( .A1(n3126), .A2(a[15]), .ZN(n3131) );
  INV_X1 U1564 ( .A(n3125), .ZN(n3126) );
  NAND2_X1 U1566 ( .A1(n3190), .A2(n3184), .ZN(n884) );
  AOI22_X1 U1567 ( .A1(n3128), .A2(n3455), .B1(n3454), .B2(a[15]), .ZN(n1200)
         );
  XOR2_X1 U1568 ( .A(n3122), .B(n3124), .Z(n2921) );
  AOI22_X1 U1569 ( .A1(n2815), .A2(n2857), .B1(n2847), .B2(n2859), .ZN(n2817)
         );
  MUX2_X2 U1571 ( .A(n3310), .B(n3311), .S(a[23]), .Z(n2575) );
  NAND2_X1 U1572 ( .A1(n3430), .A2(n3589), .ZN(n896) );
  XNOR2_X1 U1573 ( .A(n3010), .B(a[1]), .ZN(n3001) );
  NAND2_X1 U1576 ( .A1(n1377), .A2(n45), .ZN(n1049) );
  INV_X1 U1577 ( .A(n3244), .ZN(n3247) );
  INV_X1 U1578 ( .A(n2633), .ZN(n2634) );
  NOR2_X1 U1579 ( .A1(n2572), .A2(n2571), .ZN(n2632) );
  NOR2_X1 U1580 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  NOR2_X1 U1581 ( .A1(a[25]), .A2(n2145), .ZN(n2569) );
  NOR2_X1 U1586 ( .A1(n3251), .A2(n3250), .ZN(n2541) );
  NAND2_X1 U1588 ( .A1(n2479), .A2(n2480), .ZN(n2483) );
  INV_X1 U1589 ( .A(n2480), .ZN(n2482) );
  NOR2_X1 U1590 ( .A1(n2340), .A2(n2518), .ZN(n2339) );
  OAI21_X1 U1591 ( .B1(n86), .B2(n3118), .A(n2349), .ZN(n2348) );
  NOR2_X1 U1592 ( .A1(n100), .A2(b[14]), .ZN(n2909) );
  NAND2_X2 U1593 ( .A1(n1721), .A2(n58), .ZN(n2240) );
  NOR2_X1 U1594 ( .A1(n3128), .A2(n3065), .ZN(n2825) );
  NAND2_X1 U1595 ( .A1(n4045), .A2(a[8]), .ZN(n2780) );
  NAND2_X1 U1596 ( .A1(n3187), .A2(n3186), .ZN(n3188) );
  INV_X1 U1597 ( .A(n2596), .ZN(n2598) );
  INV_X1 U1598 ( .A(n2486), .ZN(n2487) );
  AOI21_X1 U1599 ( .B1(n2629), .B2(n2628), .A(n2627), .ZN(n2675) );
  NAND2_X1 U1600 ( .A1(n1209), .A2(a[11]), .ZN(n494) );
  NAND3_X1 U1601 ( .A1(n2887), .A2(n2886), .A3(n1751), .ZN(n631) );
  NOR2_X1 U1602 ( .A1(n2698), .A2(n1047), .ZN(n2699) );
  MUX2_X2 U1603 ( .A(n3120), .B(n3119), .S(n2697), .Z(n2698) );
  NAND2_X1 U1604 ( .A1(n1049), .A2(n1048), .ZN(n1047) );
  NAND2_X1 U1605 ( .A1(n4045), .A2(a[23]), .ZN(n1048) );
  INV_X1 U1606 ( .A(n2618), .ZN(n2621) );
  AOI21_X1 U1608 ( .B1(n2589), .B2(n2394), .A(n2594), .ZN(n2627) );
  AOI21_X1 U1611 ( .B1(n3113), .B2(n97), .A(n2108), .ZN(n2107) );
  NOR2_X1 U1612 ( .A1(n2109), .A2(n97), .ZN(n2108) );
  XNOR2_X1 U1614 ( .A(n2754), .B(n2753), .ZN(n2775) );
  NAND2_X1 U1615 ( .A1(n2752), .A2(n2751), .ZN(n2754) );
  INV_X1 U1616 ( .A(n2750), .ZN(n2752) );
  INV_X1 U1617 ( .A(n3221), .ZN(n3223) );
  INV_X1 U1618 ( .A(n1283), .ZN(n770) );
  INV_X1 U1619 ( .A(n2514), .ZN(n2446) );
  NOR2_X1 U1620 ( .A1(n2245), .A2(n2486), .ZN(n740) );
  NAND3_X1 U1621 ( .A1(n2473), .A2(n35), .A3(n2474), .ZN(n1157) );
  NAND2_X1 U1622 ( .A1(n2422), .A2(n2421), .ZN(n2568) );
  INV_X1 U1623 ( .A(n2508), .ZN(n2421) );
  XNOR2_X1 U1625 ( .A(n97), .B(n3498), .ZN(n2913) );
  OR2_X2 U1626 ( .A1(n1835), .A2(n3534), .ZN(n1995) );
  INV_X1 U1627 ( .A(n2861), .ZN(n2862) );
  NOR2_X1 U1628 ( .A1(n2275), .A2(n2963), .ZN(n2964) );
  NAND2_X1 U1629 ( .A1(n3409), .A2(n3200), .ZN(n640) );
  INV_X2 U1630 ( .A(n3329), .ZN(n988) );
  INV_X1 U1632 ( .A(n2105), .ZN(n2845) );
  NAND3_X1 U1634 ( .A1(n1127), .A2(n1126), .A3(n1531), .ZN(n1533) );
  INV_X2 U1637 ( .A(n76), .ZN(n1459) );
  NAND2_X1 U1638 ( .A1(n1832), .A2(n1703), .ZN(n1389) );
  NOR2_X1 U1640 ( .A1(n2705), .A2(n2704), .ZN(n2706) );
  MUX2_X1 U1641 ( .A(n3120), .B(n3119), .S(n45), .Z(n2704) );
  MUX2_X2 U1642 ( .A(n4045), .B(n1377), .S(n3589), .Z(n2705) );
  NOR2_X1 U1643 ( .A1(n2700), .A2(n2699), .ZN(n2750) );
  NAND2_X1 U1644 ( .A1(n2700), .A2(n2699), .ZN(n2751) );
  INV_X1 U1645 ( .A(n2666), .ZN(n2670) );
  AOI21_X1 U1646 ( .B1(n2628), .B2(n2629), .A(n2627), .ZN(n1348) );
  NOR2_X1 U1647 ( .A1(n2662), .A2(n2661), .ZN(n2663) );
  NOR2_X1 U1648 ( .A1(a[25]), .A2(n1651), .ZN(n2661) );
  MUX2_X1 U1649 ( .A(n2691), .B(n2692), .S(n2301), .Z(n2714) );
  NAND2_X1 U1650 ( .A1(n2688), .A2(n2613), .ZN(n2692) );
  NAND2_X1 U1651 ( .A1(n2690), .A2(a[25]), .ZN(n2691) );
  NAND2_X2 U1652 ( .A1(n1979), .A2(n3280), .ZN(n3283) );
  NAND3_X1 U1653 ( .A1(n662), .A2(n3133), .A3(n347), .ZN(n757) );
  INV_X1 U1654 ( .A(n347), .ZN(n1851) );
  INV_X1 U1655 ( .A(n1926), .ZN(n657) );
  NAND2_X1 U1656 ( .A1(n71), .A2(n1926), .ZN(n660) );
  NAND2_X1 U1660 ( .A1(n3323), .A2(n56), .ZN(n1725) );
  NAND2_X1 U1661 ( .A1(n3329), .A2(n3139), .ZN(n1724) );
  NAND2_X1 U1662 ( .A1(n155), .A2(a[7]), .ZN(n1756) );
  NOR2_X1 U1664 ( .A1(n3304), .A2(n2366), .ZN(n2365) );
  NAND2_X1 U1665 ( .A1(n3522), .A2(n3409), .ZN(n1694) );
  INV_X1 U1666 ( .A(n3384), .ZN(n3314) );
  NAND2_X2 U1667 ( .A1(n2354), .A2(n2355), .ZN(n2351) );
  NOR2_X2 U1668 ( .A1(n3306), .A2(n3073), .ZN(n2353) );
  NAND2_X1 U1669 ( .A1(n3203), .A2(a[1]), .ZN(n825) );
  NAND2_X1 U1671 ( .A1(n3119), .A2(n2045), .ZN(n700) );
  NAND2_X1 U1672 ( .A1(n3120), .A2(a[1]), .ZN(n699) );
  NAND2_X1 U1674 ( .A1(n4045), .A2(n2356), .ZN(n702) );
  MUX2_X1 U1675 ( .A(n1262), .B(n3454), .S(n205), .Z(n3315) );
  NAND2_X1 U1676 ( .A1(n3453), .A2(a[7]), .ZN(n816) );
  NOR3_X1 U1677 ( .A1(n3509), .A2(n3508), .A3(n3506), .ZN(n3507) );
  NOR2_X1 U1678 ( .A1(n3522), .A2(n3515), .ZN(n3506) );
  XNOR2_X1 U1679 ( .A(n2356), .B(n2020), .ZN(n3496) );
  INV_X1 U1680 ( .A(n3498), .ZN(n2020) );
  INV_X1 U1684 ( .A(n3368), .ZN(n690) );
  INV_X1 U1685 ( .A(n2648), .ZN(n2649) );
  INV_X1 U1686 ( .A(n2645), .ZN(n2643) );
  MUX2_X2 U1687 ( .A(n2742), .B(n3076), .S(n2613), .Z(n3592) );
  NOR2_X1 U1688 ( .A1(n3803), .A2(n3369), .ZN(n2195) );
  INV_X1 U1689 ( .A(n2734), .ZN(n2684) );
  AOI21_X1 U1690 ( .B1(n1705), .B2(n3644), .A(n3643), .ZN(n3843) );
  MUX2_X1 U1692 ( .A(n1721), .B(n3208), .S(a[25]), .Z(n3841) );
  XNOR2_X1 U1693 ( .A(n2716), .B(n2701), .ZN(n2726) );
  XNOR2_X1 U1694 ( .A(n2715), .B(n2714), .ZN(n2716) );
  OAI21_X1 U1695 ( .B1(n3377), .B2(n3374), .A(n3375), .ZN(n3575) );
  NOR2_X1 U1696 ( .A1(n2739), .A2(n2738), .ZN(n3583) );
  MUX2_X2 U1697 ( .A(n2654), .B(n2296), .S(n45), .Z(n2738) );
  MUX2_X2 U1698 ( .A(n2737), .B(n2736), .S(a[24]), .Z(n2739) );
  INV_X1 U1699 ( .A(n2731), .ZN(n2732) );
  NOR2_X1 U1700 ( .A1(n3595), .A2(n2731), .ZN(n2735) );
  INV_X1 U1701 ( .A(n3595), .ZN(n2733) );
  INV_X1 U1702 ( .A(n3096), .ZN(n3100) );
  INV_X1 U1703 ( .A(n1631), .ZN(n3271) );
  MUX2_X2 U1704 ( .A(n4085), .B(n1261), .S(n1784), .Z(n3319) );
  MUX2_X1 U1705 ( .A(n1262), .B(n3454), .S(a[7]), .Z(n3081) );
  BUF_X4 U1706 ( .A(n432), .Z(n602) );
  NAND2_X1 U1708 ( .A1(n922), .A2(a[7]), .ZN(n1034) );
  MUX2_X1 U1709 ( .A(n3513), .B(n3512), .S(n2356), .Z(n3514) );
  NAND2_X1 U1710 ( .A1(n1088), .A2(n99), .ZN(n3477) );
  MUX2_X2 U1711 ( .A(n1016), .B(n3472), .S(n3538), .Z(n3473) );
  INV_X1 U1712 ( .A(n3479), .ZN(n3543) );
  XNOR2_X1 U1713 ( .A(n3434), .B(n3433), .ZN(n3436) );
  NOR2_X1 U1714 ( .A1(n3647), .A2(n3646), .ZN(n3650) );
  NAND2_X1 U1715 ( .A1(n3647), .A2(n3646), .ZN(n3651) );
  XNOR2_X1 U1716 ( .A(n3844), .B(n3843), .ZN(n3654) );
  NOR2_X1 U1717 ( .A1(n2969), .A2(n2967), .ZN(n1182) );
  NAND2_X1 U1718 ( .A1(n987), .A2(n3362), .ZN(n1170) );
  INV_X1 U1719 ( .A(n2261), .ZN(n501) );
  NAND2_X1 U1722 ( .A1(n3434), .A2(n3433), .ZN(n3395) );
  INV_X1 U1723 ( .A(n3434), .ZN(n2182) );
  XNOR2_X1 U1724 ( .A(n2743), .B(n3595), .ZN(n3581) );
  XNOR2_X1 U1725 ( .A(n3593), .B(n3592), .ZN(n2743) );
  AOI21_X1 U1726 ( .B1(n2712), .B2(n2711), .A(n2708), .ZN(n2729) );
  INV_X1 U1727 ( .A(n2710), .ZN(n2708) );
  NAND2_X1 U1728 ( .A1(n3576), .A2(n3575), .ZN(n3711) );
  NOR2_X2 U1729 ( .A1(n62), .A2(n3829), .ZN(n2344) );
  NAND2_X1 U1730 ( .A1(n3400), .A2(n4159), .ZN(n3335) );
  NAND2_X1 U1731 ( .A1(n915), .A2(n1016), .ZN(n3552) );
  INV_X1 U1732 ( .A(n3544), .ZN(n3548) );
  NAND2_X1 U1735 ( .A1(n3654), .A2(n3648), .ZN(n3837) );
  AOI21_X1 U1736 ( .B1(n3651), .B2(n3649), .A(n3650), .ZN(n3648) );
  NAND2_X2 U1737 ( .A1(n3684), .A2(n3683), .ZN(n3917) );
  INV_X1 U1738 ( .A(n3682), .ZN(n3684) );
  NAND2_X1 U1739 ( .A1(n3917), .A2(n14), .ZN(n3916) );
  INV_X1 U1740 ( .A(n3917), .ZN(n3918) );
  INV_X1 U1741 ( .A(n3916), .ZN(n3921) );
  NOR2_X2 U1742 ( .A1(n3720), .A2(n1847), .ZN(n3620) );
  NOR2_X1 U1743 ( .A1(n3588), .A2(n3587), .ZN(n3600) );
  NOR2_X1 U1744 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  AOI21_X1 U1745 ( .B1(n3586), .B2(n3585), .A(n3584), .ZN(n3588) );
  INV_X1 U1746 ( .A(n3581), .ZN(n3586) );
  XNOR2_X1 U1747 ( .A(n3598), .B(n3647), .ZN(n3599) );
  INV_X1 U1748 ( .A(n3699), .ZN(n3700) );
  INV_X1 U1749 ( .A(n3683), .ZN(n3615) );
  INV_X2 U1750 ( .A(n931), .ZN(n873) );
  INV_X1 U1753 ( .A(n3364), .ZN(n694) );
  NOR2_X1 U1758 ( .A1(n3655), .A2(n3847), .ZN(n3668) );
  INV_X1 U1759 ( .A(n3837), .ZN(n3655) );
  INV_X1 U1760 ( .A(n3838), .ZN(n3669) );
  NOR2_X2 U1761 ( .A1(n3920), .A2(n3917), .ZN(n3928) );
  NAND2_X1 U1762 ( .A1(n3898), .A2(n3895), .ZN(n3896) );
  NAND2_X2 U1763 ( .A1(n3901), .A2(n3894), .ZN(n3984) );
  INV_X1 U1764 ( .A(n3812), .ZN(n3800) );
  INV_X1 U1767 ( .A(n4017), .ZN(n3996) );
  NAND3_X1 U1768 ( .A1(n852), .A2(n4019), .A3(n851), .ZN(n3852) );
  NOR2_X1 U1769 ( .A1(n3612), .A2(n3720), .ZN(n851) );
  INV_X1 U1770 ( .A(n4025), .ZN(n853) );
  NOR2_X2 U1771 ( .A1(n3618), .A2(n3617), .ZN(n856) );
  INV_X1 U1772 ( .A(n3658), .ZN(n3864) );
  NAND2_X1 U1773 ( .A1(n3600), .A2(n3599), .ZN(n3838) );
  INV_X1 U1774 ( .A(n3830), .ZN(n3907) );
  NOR2_X1 U1777 ( .A1(n4005), .A2(n4008), .ZN(n3739) );
  INV_X1 U1779 ( .A(n3936), .ZN(n3937) );
  AOI21_X1 U1780 ( .B1(n3869), .B2(n3868), .A(n3867), .ZN(n3880) );
  NAND3_X1 U1781 ( .A1(n3866), .A2(n3865), .A3(n3864), .ZN(n3867) );
  NAND3_X1 U1782 ( .A1(n3859), .A2(n3858), .A3(n3857), .ZN(n3860) );
  NAND2_X1 U1783 ( .A1(n3856), .A2(n3855), .ZN(n3858) );
  INV_X1 U1784 ( .A(n3853), .ZN(n3855) );
  NOR3_X1 U1785 ( .A1(n3919), .A2(n3876), .A3(n3875), .ZN(n3877) );
  INV_X1 U1786 ( .A(n3874), .ZN(n3876) );
  NAND3_X1 U1787 ( .A1(n3728), .A2(n61), .A3(n3722), .ZN(n3723) );
  INV_X1 U1788 ( .A(n3728), .ZN(n2307) );
  AOI22_X1 U1789 ( .A1(n3957), .A2(n1617), .B1(n1570), .B2(n1311), .ZN(n3958)
         );
  NAND2_X1 U1790 ( .A1(n3780), .A2(n3779), .ZN(n3782) );
  INV_X1 U1791 ( .A(n3809), .ZN(n3786) );
  NOR2_X1 U1793 ( .A1(n3815), .A2(n3814), .ZN(n3816) );
  XNOR2_X1 U1794 ( .A(n1184), .B(n3778), .ZN(\d[11] ) );
  AOI22_X1 U1795 ( .A1(n3783), .A2(n1186), .B1(n1185), .B2(n3784), .ZN(n1184)
         );
  NAND2_X1 U1796 ( .A1(n3638), .A2(n3637), .ZN(n3622) );
  NAND2_X1 U1797 ( .A1(n3864), .A2(n3838), .ZN(n3621) );
  XNOR2_X1 U1798 ( .A(n3771), .B(n3770), .ZN(\d[8]_BAR ) );
  AOI21_X1 U1799 ( .B1(n3769), .B2(n3768), .A(n3767), .ZN(n3770) );
  INV_X4 U1801 ( .A(n3265), .ZN(n2358) );
  NAND2_X1 U1803 ( .A1(n3779), .A2(n516), .ZN(n1186) );
  INV_X1 U1804 ( .A(n2476), .ZN(n737) );
  INV_X4 U1805 ( .A(a[9]), .ZN(n3139) );
  INV_X4 U1807 ( .A(n3090), .ZN(n3089) );
  INV_X4 U1809 ( .A(n3237), .ZN(n1518) );
  INV_X4 U1810 ( .A(n2038), .ZN(n2031) );
  INV_X4 U1811 ( .A(n3839), .ZN(n2109) );
  AND2_X4 U1812 ( .A1(n2315), .A2(a[11]), .ZN(n441) );
  XNOR2_X1 U1813 ( .A(n3784), .B(n3783), .ZN(n442) );
  NOR2_X2 U1814 ( .A1(n2791), .A2(n2784), .ZN(n2829) );
  XNOR2_X1 U1815 ( .A(n3498), .B(n2228), .ZN(n444) );
  AOI21_X1 U1816 ( .B1(n613), .B2(n3464), .A(n3463), .ZN(n3484) );
  INV_X4 U1818 ( .A(n2503), .ZN(n2252) );
  XOR2_X1 U1819 ( .A(a[23]), .B(n3498), .Z(n445) );
  NOR2_X1 U1821 ( .A1(n1383), .A2(n3443), .ZN(n597) );
  INV_X2 U1822 ( .A(n2858), .ZN(n2860) );
  AND2_X2 U1823 ( .A1(n3193), .A2(n3194), .ZN(n449) );
  AND2_X4 U1824 ( .A1(n922), .A2(a[24]), .ZN(n450) );
  AND2_X2 U1825 ( .A1(n2315), .A2(a[8]), .ZN(n451) );
  AND2_X2 U1826 ( .A1(n1659), .A2(n1221), .ZN(n452) );
  INV_X4 U1827 ( .A(n2847), .ZN(n2814) );
  NAND2_X2 U1828 ( .A1(n2848), .A2(n1919), .ZN(n2853) );
  AND2_X4 U1829 ( .A1(n2278), .A2(n3193), .ZN(n454) );
  INV_X4 U1830 ( .A(n3288), .ZN(n1440) );
  AND2_X4 U1832 ( .A1(n3177), .A2(n2355), .ZN(n459) );
  INV_X2 U1833 ( .A(n1541), .ZN(n743) );
  NOR2_X1 U1834 ( .A1(n2592), .A2(n2591), .ZN(n2593) );
  INV_X1 U1835 ( .A(n2593), .ZN(n2594) );
  NAND2_X1 U1836 ( .A1(n3486), .A2(n3484), .ZN(n3492) );
  INV_X1 U1837 ( .A(n3492), .ZN(n1967) );
  NOR2_X2 U1838 ( .A1(n3323), .A2(n3409), .ZN(n462) );
  INV_X1 U1839 ( .A(n3779), .ZN(n3774) );
  XNOR2_X1 U1840 ( .A(a[20]), .B(n1651), .ZN(n467) );
  INV_X1 U1841 ( .A(n4019), .ZN(n3993) );
  INV_X1 U1842 ( .A(a[11]), .ZN(n2258) );
  NAND2_X2 U1844 ( .A1(n849), .A2(n2678), .ZN(n3574) );
  AOI22_X1 U1846 ( .A1(n2483), .A2(n2158), .B1(n2481), .B2(n2482), .ZN(n2484)
         );
  NOR2_X2 U1847 ( .A1(n1120), .A2(n4050), .ZN(n3183) );
  INV_X4 U1850 ( .A(a[17]), .ZN(n1554) );
  OAI22_X1 U1851 ( .A1(n2997), .A2(n2535), .B1(n3010), .B2(n2534), .ZN(n3250)
         );
  NAND2_X1 U1852 ( .A1(n3176), .A2(n3217), .ZN(n475) );
  INV_X2 U1853 ( .A(n3538), .ZN(n916) );
  INV_X1 U1854 ( .A(n3176), .ZN(n1081) );
  INV_X1 U1856 ( .A(n2400), .ZN(n2057) );
  INV_X4 U1857 ( .A(a[22]), .ZN(n2697) );
  INV_X4 U1858 ( .A(a[15]), .ZN(n3128) );
  AOI22_X1 U1862 ( .A1(n2670), .A2(n2669), .B1(n2668), .B2(n2667), .ZN(n2671)
         );
  NAND3_X2 U1863 ( .A1(n480), .A2(n2599), .A3(n2601), .ZN(n728) );
  NOR2_X2 U1865 ( .A1(n2502), .A2(n2493), .ZN(n477) );
  NAND2_X2 U1866 ( .A1(n2253), .A2(n2252), .ZN(n478) );
  XNOR2_X2 U1867 ( .A(n479), .B(n2626), .ZN(n2599) );
  NAND2_X2 U1868 ( .A1(n1188), .A2(n2629), .ZN(n479) );
  NAND2_X2 U1870 ( .A1(n2491), .A2(n2492), .ZN(n2602) );
  INV_X8 U1872 ( .A(n482), .ZN(n3200) );
  NOR2_X2 U1873 ( .A1(n2498), .A2(n2572), .ZN(n2620) );
  NOR2_X2 U1874 ( .A1(n484), .A2(n483), .ZN(n2572) );
  AND2_X2 U1875 ( .A1(n482), .A2(n2613), .ZN(n483) );
  NAND2_X2 U1876 ( .A1(n2382), .A2(n2145), .ZN(n482) );
  NOR2_X2 U1877 ( .A1(n2613), .A2(n3453), .ZN(n484) );
  NAND2_X2 U1878 ( .A1(n2382), .A2(n2785), .ZN(n481) );
  INV_X2 U1879 ( .A(n1068), .ZN(n3045) );
  NAND2_X2 U1880 ( .A1(n1265), .A2(n2385), .ZN(n1068) );
  NAND2_X2 U1881 ( .A1(n489), .A2(n488), .ZN(n2385) );
  NAND2_X1 U1882 ( .A1(n2040), .A2(n2990), .ZN(n488) );
  NOR2_X1 U1883 ( .A1(n2991), .A2(n3026), .ZN(n491) );
  NAND2_X2 U1884 ( .A1(n1236), .A2(n2155), .ZN(n3025) );
  NOR3_X2 U1885 ( .A1(n462), .A2(n495), .A3(n2153), .ZN(n1236) );
  NOR2_X2 U1888 ( .A1(n498), .A2(n497), .ZN(n2155) );
  NAND2_X2 U1890 ( .A1(n501), .A2(n2262), .ZN(n499) );
  NAND2_X2 U1891 ( .A1(n500), .A2(n3372), .ZN(n2262) );
  NAND2_X2 U1892 ( .A1(n1384), .A2(n446), .ZN(n500) );
  NOR2_X2 U1893 ( .A1(n1384), .A2(n446), .ZN(n2261) );
  NAND2_X2 U1894 ( .A1(n1429), .A2(n1428), .ZN(n726) );
  NOR2_X2 U1895 ( .A1(n502), .A2(n3101), .ZN(n3096) );
  AOI21_X2 U1896 ( .B1(n502), .B2(n3101), .A(n68), .ZN(n2166) );
  NAND2_X2 U1897 ( .A1(n1313), .A2(n503), .ZN(n1727) );
  BUF_X4 U1899 ( .A(n1647), .Z(n505) );
  NAND2_X2 U1900 ( .A1(n1634), .A2(n1647), .ZN(n1072) );
  NAND2_X1 U1901 ( .A1(n3245), .A2(n1647), .ZN(n1842) );
  NAND3_X2 U1904 ( .A1(n1868), .A2(n1867), .A3(n1865), .ZN(n3092) );
  NAND2_X1 U1905 ( .A1(n508), .A2(n398), .ZN(n507) );
  NAND2_X2 U1906 ( .A1(n3091), .A2(n1661), .ZN(n510) );
  INV_X2 U1907 ( .A(n511), .ZN(n1805) );
  NOR2_X2 U1908 ( .A1(n3493), .A2(n1967), .ZN(n3760) );
  NOR2_X2 U1909 ( .A1(n3482), .A2(n3487), .ZN(n3493) );
  NAND2_X1 U1910 ( .A1(n1969), .A2(n3451), .ZN(n512) );
  NAND2_X2 U1911 ( .A1(n1351), .A2(n1352), .ZN(n513) );
  XNOR2_X1 U1912 ( .A(n1186), .B(n442), .ZN(\d[10]_BAR ) );
  INV_X2 U1913 ( .A(n1748), .ZN(n3452) );
  NAND2_X2 U1914 ( .A1(n518), .A2(n517), .ZN(n1748) );
  OAI21_X2 U1916 ( .B1(n830), .B2(n3050), .A(n3049), .ZN(n917) );
  NOR2_X2 U1917 ( .A1(n539), .A2(n1661), .ZN(n1711) );
  NAND2_X2 U1918 ( .A1(n1460), .A2(n1461), .ZN(n1661) );
  NAND2_X2 U1919 ( .A1(n1575), .A2(n1574), .ZN(n519) );
  NAND2_X2 U1920 ( .A1(n1298), .A2(n3050), .ZN(n3088) );
  NAND2_X2 U1921 ( .A1(n3739), .A2(n4023), .ZN(n537) );
  NOR2_X2 U1922 ( .A1(n3963), .A2(n1098), .ZN(n521) );
  OAI21_X2 U1923 ( .B1(n523), .B2(n3603), .A(n522), .ZN(n3735) );
  NOR2_X4 U1924 ( .A1(n819), .A2(n818), .ZN(n3603) );
  NOR2_X2 U1925 ( .A1(n1771), .A2(n1260), .ZN(n523) );
  NAND3_X2 U1926 ( .A1(n3070), .A2(n2193), .A3(n1890), .ZN(n524) );
  INV_X4 U1927 ( .A(n524), .ZN(n1659) );
  NAND2_X1 U1928 ( .A1(a[19]), .A2(n524), .ZN(n2940) );
  INV_X2 U1929 ( .A(n525), .ZN(n1386) );
  NOR2_X2 U1930 ( .A1(n1980), .A2(n3275), .ZN(n525) );
  NOR2_X2 U1931 ( .A1(n526), .A2(n3253), .ZN(n3275) );
  NOR2_X2 U1932 ( .A1(n540), .A2(n3254), .ZN(n526) );
  NOR2_X4 U1933 ( .A1(n2392), .A2(n3274), .ZN(n1980) );
  INV_X4 U1934 ( .A(n1695), .ZN(n2392) );
  NAND2_X2 U1935 ( .A1(n2013), .A2(n2105), .ZN(n955) );
  NAND2_X2 U1936 ( .A1(n532), .A2(n531), .ZN(n2105) );
  OAI22_X2 U1940 ( .A1(n2821), .A2(n2822), .B1(n3306), .B2(n2820), .ZN(n531)
         );
  AOI22_X2 U1941 ( .A1(n2997), .A2(n2824), .B1(n92), .B2(n2823), .ZN(n532) );
  NAND2_X2 U1942 ( .A1(n534), .A2(n533), .ZN(\d[28] ) );
  NAND2_X2 U1943 ( .A1(n535), .A2(n282), .ZN(n534) );
  NOR2_X2 U1945 ( .A1(n1482), .A2(n4015), .ZN(n536) );
  NAND2_X2 U1946 ( .A1(n537), .A2(n2381), .ZN(n3741) );
  NAND3_X1 U1947 ( .A1(n537), .A2(n3742), .A3(n2381), .ZN(n3743) );
  INV_X2 U1948 ( .A(n539), .ZN(n538) );
  NAND3_X2 U1949 ( .A1(n3932), .A2(n3930), .A3(n3931), .ZN(\d[35]_BAR ) );
  NAND3_X2 U1950 ( .A1(n1481), .A2(n2548), .A3(n2071), .ZN(n540) );
  NAND2_X2 U1951 ( .A1(n542), .A2(n1291), .ZN(n541) );
  INV_X2 U1952 ( .A(n544), .ZN(n542) );
  NAND3_X2 U1954 ( .A1(n3117), .A2(n1854), .A3(n3114), .ZN(n3221) );
  NAND2_X2 U1955 ( .A1(n3116), .A2(n3115), .ZN(n3222) );
  NAND3_X2 U1956 ( .A1(n1955), .A2(n805), .A3(n3276), .ZN(n1956) );
  INV_X4 U1959 ( .A(n3242), .ZN(n1624) );
  INV_X4 U1961 ( .A(n2004), .ZN(n2007) );
  NAND2_X2 U1962 ( .A1(n550), .A2(n549), .ZN(n2004) );
  INV_X2 U1963 ( .A(n1132), .ZN(n551) );
  INV_X2 U1964 ( .A(n553), .ZN(n552) );
  NAND2_X2 U1965 ( .A1(n2003), .A2(n3295), .ZN(n553) );
  NOR2_X2 U1966 ( .A1(n2305), .A2(n3248), .ZN(n1132) );
  NAND2_X2 U1967 ( .A1(n556), .A2(n555), .ZN(n1954) );
  INV_X4 U1968 ( .A(n1599), .ZN(n557) );
  NOR2_X4 U1969 ( .A1(n558), .A2(n557), .ZN(n3003) );
  NAND2_X2 U1970 ( .A1(n1598), .A2(n559), .ZN(n558) );
  NAND2_X2 U1971 ( .A1(n1598), .A2(n1599), .ZN(n2819) );
  NOR2_X2 U1972 ( .A1(n3329), .A2(n88), .ZN(n1181) );
  NAND2_X2 U1974 ( .A1(n996), .A2(n560), .ZN(n990) );
  INV_X4 U1975 ( .A(n2904), .ZN(n1198) );
  NAND2_X2 U1976 ( .A1(n1060), .A2(n2295), .ZN(n2904) );
  NAND2_X2 U1977 ( .A1(n562), .A2(n561), .ZN(n2295) );
  NAND2_X2 U1978 ( .A1(n625), .A2(n2051), .ZN(n561) );
  NAND2_X2 U1979 ( .A1(n1393), .A2(n2864), .ZN(n562) );
  NAND2_X2 U1980 ( .A1(n564), .A2(n563), .ZN(n1060) );
  NAND2_X2 U1981 ( .A1(n72), .A2(n1595), .ZN(n563) );
  NAND2_X2 U1983 ( .A1(n567), .A2(n565), .ZN(n3367) );
  NOR3_X2 U1984 ( .A1(n3040), .A2(n3039), .A3(n3042), .ZN(n565) );
  NOR2_X2 U1985 ( .A1(n991), .A2(n3339), .ZN(n3042) );
  NAND2_X2 U1986 ( .A1(n3015), .A2(n3014), .ZN(n3029) );
  NOR2_X2 U1987 ( .A1(n566), .A2(n3031), .ZN(n3040) );
  INV_X2 U1988 ( .A(n3030), .ZN(n566) );
  NAND2_X2 U1989 ( .A1(n3340), .A2(n3038), .ZN(n567) );
  NAND2_X2 U1990 ( .A1(n991), .A2(n3339), .ZN(n3038) );
  INV_X2 U1991 ( .A(n1931), .ZN(n570) );
  INV_X8 U1992 ( .A(n572), .ZN(n3034) );
  NAND2_X4 U1993 ( .A1(n3034), .A2(n3010), .ZN(n2980) );
  INV_X8 U1994 ( .A(n2924), .ZN(n3010) );
  OAI22_X2 U1995 ( .A1(n3644), .A2(n573), .B1(a[12]), .B2(n2980), .ZN(n1942)
         );
  INV_X1 U1996 ( .A(n2101), .ZN(n573) );
  XNOR2_X1 U1997 ( .A(n2924), .B(a[11]), .ZN(n2101) );
  INV_X1 U1998 ( .A(a[4]), .ZN(n1706) );
  NAND2_X2 U1999 ( .A1(n575), .A2(n576), .ZN(n1680) );
  NAND2_X2 U2000 ( .A1(n2859), .A2(n2847), .ZN(n575) );
  NAND2_X2 U2001 ( .A1(n577), .A2(n2814), .ZN(n576) );
  NAND2_X2 U2002 ( .A1(n579), .A2(n578), .ZN(n577) );
  INV_X2 U2003 ( .A(n443), .ZN(n578) );
  INV_X2 U2004 ( .A(n2095), .ZN(n579) );
  AOI22_X2 U2005 ( .A1(n1055), .A2(n2808), .B1(n2797), .B2(n2796), .ZN(n2847)
         );
  NOR2_X2 U2006 ( .A1(n2095), .A2(n443), .ZN(n2859) );
  NAND2_X2 U2008 ( .A1(n581), .A2(n2546), .ZN(n2530) );
  INV_X1 U2009 ( .A(n584), .ZN(n581) );
  NAND3_X2 U2010 ( .A1(n2524), .A2(n2523), .A3(n2522), .ZN(n2531) );
  NAND2_X1 U2011 ( .A1(n2407), .A2(n1449), .ZN(n582) );
  NAND2_X2 U2012 ( .A1(n923), .A2(a[19]), .ZN(n583) );
  NAND2_X2 U2013 ( .A1(n584), .A2(n80), .ZN(n2524) );
  NAND2_X2 U2014 ( .A1(n1824), .A2(n1823), .ZN(n584) );
  NAND2_X2 U2015 ( .A1(n1735), .A2(n2740), .ZN(n1361) );
  NOR2_X4 U2016 ( .A1(n585), .A2(n1600), .ZN(n1735) );
  NOR2_X4 U2017 ( .A1(b[9]), .A2(b[10]), .ZN(n1600) );
  AOI21_X2 U2018 ( .B1(n586), .B2(n3043), .A(n3048), .ZN(n1222) );
  NAND2_X2 U2019 ( .A1(n588), .A2(n587), .ZN(n709) );
  NAND2_X2 U2020 ( .A1(n871), .A2(n3366), .ZN(n3043) );
  INV_X2 U2021 ( .A(n3047), .ZN(n586) );
  NOR2_X2 U2022 ( .A1(n588), .A2(n587), .ZN(n3047) );
  NAND2_X2 U2023 ( .A1(n869), .A2(n868), .ZN(n587) );
  NOR2_X2 U2026 ( .A1(n735), .A2(n733), .ZN(n2245) );
  AOI21_X2 U2027 ( .B1(n735), .B2(n733), .A(n1567), .ZN(n2246) );
  NOR2_X2 U2028 ( .A1(n1657), .A2(n3781), .ZN(n663) );
  NAND2_X2 U2029 ( .A1(n591), .A2(n589), .ZN(n1657) );
  NAND3_X2 U2030 ( .A1(n590), .A2(n596), .A3(n593), .ZN(n589) );
  OAI21_X1 U2031 ( .B1(n597), .B2(n592), .A(n3444), .ZN(n591) );
  INV_X1 U2032 ( .A(n593), .ZN(n592) );
  AOI22_X2 U2033 ( .A1(n1551), .A2(n1552), .B1(n4143), .B2(n3418), .ZN(n598)
         );
  OAI21_X2 U2034 ( .B1(n595), .B2(n594), .A(n3443), .ZN(n593) );
  INV_X2 U2036 ( .A(n597), .ZN(n596) );
  NOR2_X2 U2037 ( .A1(n3417), .A2(n3416), .ZN(n3443) );
  INV_X2 U2038 ( .A(n3420), .ZN(n3397) );
  NAND2_X2 U2040 ( .A1(n600), .A2(n1172), .ZN(n1019) );
  NAND2_X2 U2041 ( .A1(n985), .A2(n1214), .ZN(n600) );
  NAND2_X2 U2042 ( .A1(n3538), .A2(n601), .ZN(n3465) );
  NAND2_X2 U2043 ( .A1(n604), .A2(n603), .ZN(n1485) );
  NAND2_X2 U2045 ( .A1(n606), .A2(n605), .ZN(n2404) );
  NAND2_X1 U2046 ( .A1(n2432), .A2(n2433), .ZN(n605) );
  NAND2_X2 U2047 ( .A1(n734), .A2(n1567), .ZN(n606) );
  NAND2_X2 U2048 ( .A1(n1663), .A2(n3542), .ZN(n1679) );
  AOI21_X2 U2049 ( .B1(n1396), .B2(n3545), .A(n3543), .ZN(n3542) );
  NOR2_X2 U2050 ( .A1(n1396), .A2(n3545), .ZN(n3555) );
  INV_X4 U2052 ( .A(n609), .ZN(n1908) );
  NAND2_X2 U2053 ( .A1(n611), .A2(n610), .ZN(n1911) );
  INV_X1 U2055 ( .A(n3338), .ZN(n3322) );
  INV_X2 U2056 ( .A(n3383), .ZN(n1796) );
  NOR2_X2 U2057 ( .A1(n3464), .A2(n613), .ZN(n3463) );
  NAND2_X2 U2059 ( .A1(n616), .A2(n614), .ZN(n3184) );
  AOI21_X2 U2060 ( .B1(n1231), .B2(a[10]), .A(n615), .ZN(n614) );
  NAND2_X2 U2061 ( .A1(n1493), .A2(n1494), .ZN(n616) );
  NAND2_X2 U2062 ( .A1(n2952), .A2(n1362), .ZN(n3193) );
  NOR3_X2 U2063 ( .A1(n3137), .A2(n3146), .A3(n3136), .ZN(n2952) );
  NAND2_X2 U2064 ( .A1(n620), .A2(n618), .ZN(n971) );
  NOR2_X2 U2067 ( .A1(n658), .A2(n659), .ZN(n619) );
  NAND2_X2 U2068 ( .A1(n2966), .A2(n1926), .ZN(n1173) );
  NAND2_X2 U2070 ( .A1(n622), .A2(n3302), .ZN(n1512) );
  OAI21_X1 U2071 ( .B1(n3513), .B2(a[8]), .A(n623), .ZN(n3415) );
  NAND2_X1 U2072 ( .A1(n1235), .A2(a[8]), .ZN(n623) );
  INV_X2 U2073 ( .A(n624), .ZN(n1378) );
  NAND2_X2 U2074 ( .A1(n1242), .A2(n1241), .ZN(n624) );
  INV_X2 U2075 ( .A(n2864), .ZN(n625) );
  INV_X2 U2076 ( .A(n626), .ZN(n2876) );
  NAND2_X2 U2077 ( .A1(n628), .A2(n627), .ZN(n2875) );
  NAND2_X2 U2078 ( .A1(n957), .A2(n2829), .ZN(n628) );
  AOI22_X2 U2081 ( .A1(n1444), .A2(n714), .B1(n3387), .B2(n3386), .ZN(n2368)
         );
  NOR2_X2 U2082 ( .A1(n634), .A2(n633), .ZN(n3442) );
  NOR2_X2 U2083 ( .A1(n3397), .A2(n3418), .ZN(n633) );
  NOR2_X1 U2084 ( .A1(n3396), .A2(n4143), .ZN(n634) );
  NAND2_X2 U2085 ( .A1(n635), .A2(n2794), .ZN(n2858) );
  NAND2_X2 U2086 ( .A1(n636), .A2(n2792), .ZN(n635) );
  INV_X2 U2087 ( .A(n2160), .ZN(n1403) );
  NAND2_X2 U2088 ( .A1(n2566), .A2(n2567), .ZN(n2160) );
  NAND2_X2 U2089 ( .A1(n2102), .A2(n932), .ZN(n2567) );
  NAND2_X2 U2090 ( .A1(n638), .A2(n637), .ZN(n2566) );
  INV_X2 U2091 ( .A(n932), .ZN(n637) );
  INV_X2 U2092 ( .A(n2102), .ZN(n638) );
  NAND2_X1 U2093 ( .A1(n1266), .A2(n205), .ZN(n1693) );
  NOR2_X1 U2094 ( .A1(n3958), .A2(n641), .ZN(n3959) );
  NOR3_X4 U2095 ( .A1(n1938), .A2(n4010), .A3(n1305), .ZN(n641) );
  INV_X2 U2096 ( .A(n1368), .ZN(n1204) );
  NAND2_X2 U2097 ( .A1(n23), .A2(n642), .ZN(n1368) );
  AOI21_X2 U2099 ( .B1(n644), .B2(n3228), .A(n3227), .ZN(n3265) );
  NAND2_X4 U2101 ( .A1(n645), .A2(n3194), .ZN(n3192) );
  NAND2_X1 U2102 ( .A1(n884), .A2(n645), .ZN(n883) );
  INV_X2 U2103 ( .A(n835), .ZN(n836) );
  NAND3_X2 U2104 ( .A1(n648), .A2(n647), .A3(n646), .ZN(\d[23] ) );
  NAND2_X2 U2105 ( .A1(n3914), .A2(n835), .ZN(n646) );
  INV_X2 U2106 ( .A(n649), .ZN(n648) );
  NOR2_X2 U2107 ( .A1(n835), .A2(n457), .ZN(n649) );
  OAI21_X2 U2108 ( .B1(n2068), .B2(n2069), .A(n3265), .ZN(n650) );
  NAND2_X2 U2109 ( .A1(n652), .A2(n651), .ZN(n2288) );
  NAND3_X2 U2110 ( .A1(n1299), .A2(n4151), .A3(n655), .ZN(n651) );
  NAND2_X2 U2111 ( .A1(n654), .A2(n653), .ZN(n652) );
  NAND2_X2 U2114 ( .A1(n3174), .A2(n3173), .ZN(n655) );
  AOI22_X2 U2115 ( .A1(n660), .A2(n1569), .B1(n2966), .B2(n657), .ZN(n3108) );
  AOI21_X2 U2116 ( .B1(n18), .B2(n1230), .A(n2190), .ZN(n658) );
  NOR2_X2 U2117 ( .A1(n2960), .A2(n2189), .ZN(n659) );
  NAND2_X2 U2118 ( .A1(n3788), .A2(n3787), .ZN(n3799) );
  NAND2_X2 U2119 ( .A1(n1535), .A2(n1536), .ZN(n3787) );
  NAND2_X2 U2120 ( .A1(n3806), .A2(n3803), .ZN(n3785) );
  AOI21_X2 U2121 ( .B1(n695), .B2(n694), .A(n692), .ZN(n3370) );
  NOR2_X2 U2122 ( .A1(n3776), .A2(n3783), .ZN(n664) );
  INV_X2 U2123 ( .A(n1764), .ZN(n665) );
  AOI22_X2 U2126 ( .A1(n1209), .A2(a[19]), .B1(n1863), .B2(n2407), .ZN(n667)
         );
  AOI22_X2 U2128 ( .A1(n2919), .A2(n670), .B1(n2918), .B2(n2917), .ZN(n1926)
         );
  NOR2_X4 U2129 ( .A1(n1960), .A2(n438), .ZN(n2919) );
  NAND2_X2 U2130 ( .A1(n2903), .A2(n504), .ZN(n671) );
  NAND2_X2 U2131 ( .A1(n673), .A2(n2854), .ZN(n672) );
  NAND2_X2 U2132 ( .A1(n1638), .A2(n674), .ZN(n1637) );
  NAND2_X2 U2133 ( .A1(n1594), .A2(n1593), .ZN(n674) );
  NOR2_X4 U2135 ( .A1(n2983), .A2(n3176), .ZN(n922) );
  INV_X2 U2136 ( .A(n1621), .ZN(n4012) );
  NAND3_X2 U2137 ( .A1(n1639), .A2(n1620), .A3(n1619), .ZN(n679) );
  NAND2_X2 U2138 ( .A1(n3735), .A2(n3734), .ZN(n4015) );
  NOR2_X2 U2141 ( .A1(n681), .A2(n680), .ZN(n3107) );
  AOI21_X1 U2142 ( .B1(n2234), .B2(n2233), .A(n2231), .ZN(n680) );
  NAND2_X2 U2143 ( .A1(n683), .A2(n682), .ZN(n2232) );
  INV_X2 U2144 ( .A(n2231), .ZN(n682) );
  NAND2_X2 U2145 ( .A1(n2234), .A2(n2233), .ZN(n683) );
  OAI21_X2 U2146 ( .B1(n3108), .B2(n760), .A(n759), .ZN(n1655) );
  BUF_X4 U2147 ( .A(n1655), .Z(n684) );
  NOR2_X2 U2148 ( .A1(n1655), .A2(n3229), .ZN(n756) );
  NAND2_X1 U2149 ( .A1(n1655), .A2(n3229), .ZN(n1419) );
  NAND2_X1 U2153 ( .A1(n686), .A2(n1483), .ZN(n716) );
  NAND2_X2 U2154 ( .A1(n378), .A2(n377), .ZN(n686) );
  XNOR2_X2 U2155 ( .A(n2983), .B(n2077), .ZN(n689) );
  NAND2_X2 U2157 ( .A1(n3366), .A2(n3367), .ZN(n691) );
  NOR2_X2 U2159 ( .A1(n693), .A2(n3365), .ZN(n692) );
  NAND2_X2 U2160 ( .A1(n3364), .A2(n3363), .ZN(n693) );
  NAND2_X2 U2161 ( .A1(n696), .A2(n3363), .ZN(n695) );
  INV_X2 U2162 ( .A(n3365), .ZN(n696) );
  NAND2_X2 U2163 ( .A1(n3342), .A2(n697), .ZN(n3344) );
  OAI21_X2 U2164 ( .B1(n3033), .B2(n3032), .A(n4063), .ZN(n697) );
  NAND2_X2 U2165 ( .A1(n701), .A2(n698), .ZN(n3342) );
  NOR2_X2 U2166 ( .A1(n4063), .A2(n3032), .ZN(n698) );
  NAND2_X2 U2167 ( .A1(n700), .A2(n699), .ZN(n3032) );
  INV_X2 U2168 ( .A(n3033), .ZN(n701) );
  NAND3_X1 U2169 ( .A1(n4023), .A2(n3986), .A3(n472), .ZN(n1808) );
  NOR2_X2 U2170 ( .A1(n3954), .A2(n22), .ZN(n3987) );
  NAND2_X2 U2171 ( .A1(n1703), .A2(n1832), .ZN(n1702) );
  NAND2_X2 U2172 ( .A1(n2386), .A2(n2891), .ZN(n2977) );
  INV_X4 U2174 ( .A(n3174), .ZN(n705) );
  NAND2_X2 U2175 ( .A1(n708), .A2(n706), .ZN(n1384) );
  NOR2_X2 U2177 ( .A1(n3043), .A2(n3047), .ZN(n707) );
  OAI21_X1 U2178 ( .B1(n3048), .B2(n3047), .A(n3043), .ZN(n708) );
  INV_X2 U2179 ( .A(n2934), .ZN(n2946) );
  OAI21_X2 U2181 ( .B1(n712), .B2(n714), .A(n715), .ZN(n1643) );
  NAND2_X2 U2182 ( .A1(n713), .A2(n711), .ZN(n3354) );
  INV_X2 U2183 ( .A(n712), .ZN(n711) );
  NOR2_X2 U2184 ( .A1(n1061), .A2(n3385), .ZN(n712) );
  NAND2_X2 U2185 ( .A1(n714), .A2(n715), .ZN(n713) );
  NAND2_X2 U2186 ( .A1(n1061), .A2(n3385), .ZN(n715) );
  NOR2_X1 U2188 ( .A1(n3423), .A2(n721), .ZN(n3416) );
  AOI21_X1 U2189 ( .B1(n3423), .B2(n721), .A(n3422), .ZN(n3417) );
  XNOR2_X2 U2190 ( .A(n721), .B(n3422), .ZN(n3424) );
  NAND2_X2 U2191 ( .A1(n2208), .A2(n2207), .ZN(n2159) );
  NAND2_X2 U2192 ( .A1(n722), .A2(n4158), .ZN(n2207) );
  NAND3_X2 U2193 ( .A1(n723), .A2(n1075), .A3(n4142), .ZN(n2208) );
  OAI21_X2 U2195 ( .B1(n3045), .B2(n3044), .A(n2345), .ZN(n1065) );
  NAND2_X2 U2196 ( .A1(n727), .A2(n2652), .ZN(n729) );
  NAND2_X2 U2197 ( .A1(n1269), .A2(n1268), .ZN(n2652) );
  NAND3_X2 U2198 ( .A1(n63), .A2(n2653), .A3(n728), .ZN(n730) );
  INV_X2 U2200 ( .A(n2432), .ZN(n734) );
  NOR2_X2 U2202 ( .A1(n2246), .A2(n2245), .ZN(n2489) );
  NAND2_X1 U2203 ( .A1(n2476), .A2(n1898), .ZN(n736) );
  NOR2_X2 U2204 ( .A1(n2313), .A2(n2402), .ZN(n2432) );
  INV_X2 U2205 ( .A(n2515), .ZN(n742) );
  NAND3_X2 U2206 ( .A1(n2500), .A2(n2309), .A3(n2501), .ZN(n746) );
  NOR2_X2 U2209 ( .A1(n3070), .A2(n456), .ZN(n750) );
  NOR2_X2 U2210 ( .A1(n2556), .A2(n3066), .ZN(n748) );
  NAND3_X2 U2211 ( .A1(n3266), .A2(n2358), .A3(n194), .ZN(n1882) );
  NAND2_X2 U2212 ( .A1(n753), .A2(n752), .ZN(n3571) );
  NAND2_X2 U2213 ( .A1(n1584), .A2(n1583), .ZN(n753) );
  INV_X2 U2217 ( .A(n756), .ZN(n1420) );
  NAND2_X2 U2218 ( .A1(n758), .A2(n757), .ZN(n3229) );
  NAND2_X2 U2219 ( .A1(n1785), .A2(n1851), .ZN(n758) );
  NAND2_X2 U2220 ( .A1(n3107), .A2(n3106), .ZN(n759) );
  NOR2_X2 U2221 ( .A1(n3107), .A2(n3106), .ZN(n760) );
  NAND2_X1 U2224 ( .A1(n2252), .A2(n1873), .ZN(n762) );
  NAND2_X2 U2225 ( .A1(n1355), .A2(n1356), .ZN(n764) );
  NAND3_X2 U2227 ( .A1(n767), .A2(n766), .A3(n765), .ZN(n3297) );
  NAND2_X2 U2228 ( .A1(n885), .A2(n358), .ZN(n765) );
  NAND2_X2 U2230 ( .A1(n770), .A2(n358), .ZN(n767) );
  NAND2_X2 U2231 ( .A1(n1640), .A2(n3295), .ZN(n768) );
  NAND2_X2 U2232 ( .A1(n831), .A2(n1554), .ZN(n1952) );
  OAI21_X2 U2235 ( .B1(n2242), .B2(n441), .A(n2918), .ZN(n776) );
  NAND2_X2 U2237 ( .A1(n780), .A2(n778), .ZN(n2485) );
  NAND3_X2 U2238 ( .A1(n779), .A2(n1405), .A3(n1406), .ZN(n778) );
  NAND2_X2 U2240 ( .A1(n781), .A2(n82), .ZN(n780) );
  NAND3_X2 U2241 ( .A1(n1405), .A2(n3495), .A3(n1406), .ZN(n781) );
  NOR2_X4 U2242 ( .A1(n1862), .A2(n1209), .ZN(n3535) );
  INV_X2 U2243 ( .A(n2606), .ZN(n1134) );
  NAND2_X2 U2245 ( .A1(n2309), .A2(n2501), .ZN(n940) );
  NAND2_X2 U2246 ( .A1(n782), .A2(n941), .ZN(n2605) );
  NAND2_X2 U2247 ( .A1(n1136), .A2(n2580), .ZN(n941) );
  NOR2_X4 U2248 ( .A1(n783), .A2(n2249), .ZN(n2606) );
  INV_X4 U2249 ( .A(n784), .ZN(n783) );
  NAND3_X2 U2250 ( .A1(n2601), .A2(n2602), .A3(n2250), .ZN(n784) );
  AOI22_X2 U2254 ( .A1(n81), .A2(n3462), .B1(n3466), .B2(n3465), .ZN(n3486) );
  NAND2_X2 U2255 ( .A1(n2650), .A2(n2648), .ZN(n2584) );
  NAND2_X2 U2256 ( .A1(n788), .A2(n786), .ZN(n2650) );
  INV_X2 U2257 ( .A(n787), .ZN(n786) );
  NAND2_X2 U2258 ( .A1(n1491), .A2(n1490), .ZN(n789) );
  NAND2_X2 U2260 ( .A1(n1139), .A2(n2197), .ZN(n791) );
  NAND2_X4 U2261 ( .A1(n792), .A2(n2903), .ZN(n1139) );
  NAND2_X2 U2262 ( .A1(n797), .A2(n794), .ZN(n3244) );
  NAND2_X2 U2264 ( .A1(n1377), .A2(n3016), .ZN(n796) );
  NAND2_X2 U2267 ( .A1(n831), .A2(n37), .ZN(n798) );
  NAND2_X2 U2268 ( .A1(n801), .A2(n800), .ZN(n2136) );
  NAND2_X2 U2269 ( .A1(n802), .A2(n803), .ZN(n800) );
  INV_X2 U2270 ( .A(n804), .ZN(n801) );
  NOR2_X2 U2271 ( .A1(n4054), .A2(n1166), .ZN(n804) );
  NAND3_X1 U2272 ( .A1(n1125), .A2(n3279), .A3(n805), .ZN(n1979) );
  INV_X2 U2273 ( .A(n3240), .ZN(n805) );
  AOI22_X2 U2274 ( .A1(n4204), .A2(n1282), .B1(n806), .B2(n3243), .ZN(n3248)
         );
  INV_X2 U2276 ( .A(n505), .ZN(n806) );
  NAND2_X2 U2278 ( .A1(n810), .A2(n809), .ZN(n3611) );
  NAND3_X1 U2279 ( .A1(n810), .A2(n809), .A3(n3610), .ZN(n4025) );
  AOI21_X2 U2280 ( .B1(n63), .B2(n728), .A(n893), .ZN(n3610) );
  NAND2_X2 U2283 ( .A1(n1451), .A2(n1450), .ZN(n811) );
  NAND2_X2 U2284 ( .A1(n812), .A2(n3262), .ZN(n1450) );
  INV_X2 U2285 ( .A(n1838), .ZN(n812) );
  NAND2_X2 U2286 ( .A1(n813), .A2(n1838), .ZN(n1451) );
  INV_X2 U2287 ( .A(n3262), .ZN(n813) );
  NAND3_X2 U2288 ( .A1(n453), .A2(n1130), .A3(n1129), .ZN(n3262) );
  NAND3_X2 U2289 ( .A1(n2589), .A2(n2594), .A3(n2394), .ZN(n2629) );
  NAND2_X2 U2290 ( .A1(n53), .A2(n814), .ZN(n2394) );
  INV_X2 U2291 ( .A(n2588), .ZN(n814) );
  NAND2_X2 U2292 ( .A1(n2587), .A2(n2586), .ZN(n2589) );
  INV_X2 U2294 ( .A(n87), .ZN(n1976) );
  NAND2_X2 U2295 ( .A1(n436), .A2(n3316), .ZN(n3351) );
  NOR2_X2 U2296 ( .A1(n3315), .A2(n815), .ZN(n3316) );
  OAI21_X1 U2297 ( .B1(n87), .B2(a[7]), .A(n816), .ZN(n815) );
  NAND3_X1 U2298 ( .A1(n3070), .A2(n474), .A3(n2193), .ZN(n3071) );
  INV_X1 U2299 ( .A(n3603), .ZN(n820) );
  INV_X2 U2300 ( .A(n2012), .ZN(n3749) );
  NOR2_X2 U2301 ( .A1(n829), .A2(n2261), .ZN(n828) );
  AOI22_X2 U2303 ( .A1(n3053), .A2(n1728), .B1(n83), .B2(n3052), .ZN(n830) );
  NAND2_X2 U2304 ( .A1(n831), .A2(n2613), .ZN(n2615) );
  NAND2_X2 U2305 ( .A1(n831), .A2(n95), .ZN(n2184) );
  NAND2_X2 U2307 ( .A1(n831), .A2(n54), .ZN(n1481) );
  INV_X2 U2311 ( .A(n4015), .ZN(n835) );
  OAI21_X2 U2313 ( .B1(n1878), .B2(n1492), .A(n3381), .ZN(n3577) );
  NOR2_X2 U2314 ( .A1(n839), .A2(n2671), .ZN(n1492) );
  NAND2_X2 U2315 ( .A1(n841), .A2(n840), .ZN(n839) );
  NAND3_X1 U2318 ( .A1(n75), .A2(n2655), .A3(n842), .ZN(n845) );
  NAND2_X2 U2319 ( .A1(n2615), .A2(n2614), .ZN(n843) );
  NAND2_X2 U2320 ( .A1(n2612), .A2(n2611), .ZN(n2655) );
  NAND2_X2 U2322 ( .A1(n2615), .A2(n2614), .ZN(n2664) );
  OAI21_X2 U2324 ( .B1(n2656), .B2(n848), .A(n2722), .ZN(n844) );
  NAND2_X2 U2325 ( .A1(n2646), .A2(n2645), .ZN(n2678) );
  NAND2_X2 U2326 ( .A1(n1434), .A2(n1435), .ZN(n2646) );
  NAND2_X2 U2327 ( .A1(n2677), .A2(n850), .ZN(n849) );
  NAND2_X4 U2328 ( .A1(n2644), .A2(n2643), .ZN(n2677) );
  NOR2_X1 U2329 ( .A1(n853), .A2(n3617), .ZN(n852) );
  INV_X4 U2331 ( .A(n3612), .ZN(n3722) );
  XNOR2_X2 U2333 ( .A(n3023), .B(n3024), .ZN(n1709) );
  NAND2_X2 U2334 ( .A1(n861), .A2(n858), .ZN(n3024) );
  NOR3_X2 U2337 ( .A1(n4039), .A2(n864), .A3(n862), .ZN(n3023) );
  INV_X2 U2338 ( .A(n863), .ZN(n862) );
  NAND2_X2 U2339 ( .A1(n1261), .A2(a[7]), .ZN(n863) );
  NOR2_X1 U2340 ( .A1(n3017), .A2(n432), .ZN(n864) );
  AOI22_X2 U2342 ( .A1(n3369), .A2(n3370), .B1(n1644), .B2(n867), .ZN(n3558)
         );
  INV_X4 U2343 ( .A(n3559), .ZN(n867) );
  XNOR2_X2 U2344 ( .A(n3359), .B(n3358), .ZN(n3559) );
  NAND2_X1 U2345 ( .A1(n1709), .A2(n4178), .ZN(n868) );
  NAND2_X2 U2346 ( .A1(n1030), .A2(n77), .ZN(n869) );
  NAND2_X2 U2347 ( .A1(n3367), .A2(n3368), .ZN(n871) );
  OAI22_X2 U2348 ( .A1(n960), .A2(n1705), .B1(n959), .B2(n958), .ZN(n872) );
  NAND2_X2 U2350 ( .A1(n3936), .A2(n873), .ZN(n3934) );
  NAND2_X2 U2351 ( .A1(n1892), .A2(n1999), .ZN(n3936) );
  OAI21_X2 U2352 ( .B1(n2900), .B2(n2899), .A(n89), .ZN(n875) );
  NAND2_X2 U2353 ( .A1(n878), .A2(n877), .ZN(n876) );
  INV_X2 U2354 ( .A(n2900), .ZN(n878) );
  NAND2_X2 U2355 ( .A1(n3453), .A2(a[17]), .ZN(n880) );
  NAND2_X2 U2356 ( .A1(n3200), .A2(n1554), .ZN(n881) );
  AOI22_X2 U2357 ( .A1(n882), .A2(n449), .B1(n3193), .B2(n3191), .ZN(n2042) );
  NOR2_X2 U2358 ( .A1(n3190), .A2(n3184), .ZN(n3191) );
  INV_X2 U2359 ( .A(n883), .ZN(n882) );
  INV_X4 U2360 ( .A(n3159), .ZN(n3190) );
  NAND2_X2 U2363 ( .A1(n887), .A2(n886), .ZN(n3292) );
  NAND2_X2 U2364 ( .A1(n1739), .A2(n2547), .ZN(n886) );
  NAND2_X2 U2366 ( .A1(n889), .A2(n888), .ZN(n3894) );
  NAND2_X2 U2367 ( .A1(n3888), .A2(n890), .ZN(n888) );
  NOR2_X2 U2369 ( .A1(n3892), .A2(n3963), .ZN(n3893) );
  AOI21_X2 U2370 ( .B1(n2677), .B2(n2678), .A(n2676), .ZN(n892) );
  INV_X2 U2372 ( .A(n3340), .ZN(n1963) );
  INV_X2 U2373 ( .A(n1964), .ZN(n894) );
  NAND2_X2 U2374 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X2 U2375 ( .A1(n903), .A2(n897), .ZN(n2975) );
  NOR2_X2 U2377 ( .A1(n901), .A2(n1293), .ZN(n900) );
  NAND2_X2 U2378 ( .A1(n905), .A2(n904), .ZN(n903) );
  NAND2_X1 U2379 ( .A1(n2047), .A2(n2881), .ZN(n904) );
  NAND2_X2 U2380 ( .A1(n1325), .A2(n1326), .ZN(n905) );
  NOR2_X4 U2381 ( .A1(n907), .A2(n906), .ZN(n2992) );
  NOR2_X2 U2382 ( .A1(n908), .A2(n4077), .ZN(n906) );
  AOI21_X2 U2383 ( .B1(n908), .B2(n4077), .A(n790), .ZN(n907) );
  NAND2_X2 U2385 ( .A1(n1139), .A2(n2197), .ZN(n908) );
  NAND2_X1 U2389 ( .A1(n1976), .A2(n916), .ZN(n915) );
  MUX2_X2 U2390 ( .A(n87), .B(n1121), .S(a[1]), .Z(n3474) );
  INV_X2 U2391 ( .A(n1456), .ZN(n2984) );
  INV_X2 U2392 ( .A(n1703), .ZN(n2891) );
  NAND2_X2 U2393 ( .A1(n918), .A2(n2921), .ZN(n1201) );
  NAND2_X2 U2394 ( .A1(n918), .A2(n2788), .ZN(n1107) );
  INV_X4 U2395 ( .A(n2441), .ZN(n918) );
  NAND3_X2 U2396 ( .A1(n920), .A2(n919), .A3(n1742), .ZN(n1740) );
  INV_X4 U2397 ( .A(n3108), .ZN(n919) );
  INV_X2 U2398 ( .A(n921), .ZN(n920) );
  NAND2_X2 U2399 ( .A1(n1008), .A2(n1007), .ZN(n921) );
  INV_X4 U2400 ( .A(n922), .ZN(n3512) );
  NAND2_X2 U2401 ( .A1(n922), .A2(n93), .ZN(n1765) );
  NAND2_X2 U2402 ( .A1(n923), .A2(a[15]), .ZN(n2266) );
  AOI22_X2 U2403 ( .A1(n3534), .A2(n2201), .B1(n923), .B2(a[3]), .ZN(n3401) );
  INV_X4 U2404 ( .A(n2070), .ZN(n923) );
  INV_X4 U2405 ( .A(n67), .ZN(n924) );
  NAND2_X2 U2406 ( .A1(n1204), .A2(n2321), .ZN(n925) );
  NAND2_X2 U2407 ( .A1(n1368), .A2(n1369), .ZN(n926) );
  NOR3_X2 U2409 ( .A1(n3161), .A2(n3160), .A3(n927), .ZN(n3163) );
  NOR2_X2 U2410 ( .A1(n2959), .A2(n2958), .ZN(n927) );
  INV_X4 U2412 ( .A(n928), .ZN(n3270) );
  NAND2_X2 U2413 ( .A1(n437), .A2(n2560), .ZN(n928) );
  NAND2_X2 U2414 ( .A1(n930), .A2(n929), .ZN(n2561) );
  NAND2_X2 U2415 ( .A1(n2533), .A2(n2532), .ZN(n929) );
  NOR2_X1 U2416 ( .A1(n3989), .A2(n931), .ZN(n4017) );
  NOR2_X1 U2417 ( .A1(n3953), .A2(n931), .ZN(n3960) );
  INV_X1 U2420 ( .A(n3267), .ZN(n933) );
  NOR2_X2 U2421 ( .A1(n2331), .A2(n3268), .ZN(n934) );
  NOR2_X2 U2422 ( .A1(n936), .A2(n935), .ZN(n2331) );
  NAND2_X2 U2423 ( .A1(n1307), .A2(n1308), .ZN(n938) );
  NAND2_X2 U2424 ( .A1(n2521), .A2(n2202), .ZN(n937) );
  NAND3_X2 U2425 ( .A1(n2525), .A2(n937), .A3(n938), .ZN(n1500) );
  NAND3_X2 U2427 ( .A1(n939), .A2(n941), .A3(n940), .ZN(n1373) );
  NOR2_X2 U2428 ( .A1(n2582), .A2(n943), .ZN(n942) );
  NAND2_X2 U2429 ( .A1(n2583), .A2(n2251), .ZN(n943) );
  INV_X2 U2430 ( .A(n944), .ZN(n1431) );
  NOR2_X2 U2431 ( .A1(n2158), .A2(n2481), .ZN(n944) );
  NOR2_X2 U2432 ( .A1(n948), .A2(n945), .ZN(n2481) );
  NAND2_X2 U2433 ( .A1(n947), .A2(n946), .ZN(n945) );
  AOI22_X2 U2434 ( .A1(n92), .A2(n950), .B1(n949), .B2(n2997), .ZN(n2158) );
  NAND2_X2 U2435 ( .A1(n2076), .A2(n2075), .ZN(n949) );
  INV_X4 U2441 ( .A(n2384), .ZN(n3303) );
  AOI21_X2 U2442 ( .B1(n58), .B2(n3177), .A(n1837), .ZN(n958) );
  XNOR2_X2 U2443 ( .A(n2906), .B(n3010), .ZN(n960) );
  NAND2_X1 U2444 ( .A1(n1554), .A2(n2384), .ZN(n961) );
  NAND3_X2 U2445 ( .A1(n1339), .A2(n1338), .A3(n57), .ZN(n962) );
  NAND3_X1 U2446 ( .A1(n1657), .A2(n3776), .A3(n3781), .ZN(n3446) );
  NAND2_X2 U2447 ( .A1(n963), .A2(n966), .ZN(n3776) );
  NAND2_X2 U2448 ( .A1(n70), .A2(n2368), .ZN(n964) );
  NAND2_X2 U2449 ( .A1(n1233), .A2(n1234), .ZN(n965) );
  NAND2_X2 U2450 ( .A1(n968), .A2(n967), .ZN(n966) );
  NAND2_X2 U2451 ( .A1(n1446), .A2(n1445), .ZN(n968) );
  XOR2_X1 U2452 ( .A(n559), .B(n2228), .Z(n2820) );
  NOR2_X1 U2453 ( .A1(n1449), .A2(n93), .ZN(n2214) );
  NAND2_X2 U2455 ( .A1(n971), .A2(n970), .ZN(n2968) );
  NOR2_X4 U2457 ( .A1(n1300), .A2(n2947), .ZN(n2948) );
  NAND2_X2 U2458 ( .A1(n1840), .A2(n1839), .ZN(n973) );
  NAND2_X2 U2459 ( .A1(n975), .A2(n974), .ZN(n3174) );
  NAND3_X1 U2460 ( .A1(n3170), .A2(n3171), .A3(n2317), .ZN(n974) );
  AOI21_X2 U2465 ( .B1(n2947), .B2(n1300), .A(n2946), .ZN(n977) );
  OAI22_X2 U2466 ( .A1(n2084), .A2(n3016), .B1(n3328), .B2(a[12]), .ZN(n982)
         );
  INV_X4 U2467 ( .A(n1835), .ZN(n3208) );
  NAND2_X2 U2468 ( .A1(n978), .A2(n1162), .ZN(n1211) );
  NAND2_X2 U2469 ( .A1(n980), .A2(n979), .ZN(n1162) );
  INV_X2 U2470 ( .A(n3135), .ZN(n978) );
  NOR2_X2 U2471 ( .A1(n980), .A2(n979), .ZN(n3135) );
  NAND2_X2 U2472 ( .A1(n983), .A2(n981), .ZN(n980) );
  NAND2_X2 U2474 ( .A1(n3371), .A2(n2088), .ZN(n1172) );
  INV_X2 U2475 ( .A(n2088), .ZN(n985) );
  OAI21_X2 U2476 ( .B1(n3365), .B2(n3364), .A(n3363), .ZN(n2088) );
  AOI21_X2 U2477 ( .B1(n3351), .B2(n3350), .A(n4206), .ZN(n3364) );
  NAND2_X2 U2478 ( .A1(n986), .A2(n1427), .ZN(n1171) );
  INV_X2 U2479 ( .A(n987), .ZN(n986) );
  NAND2_X2 U2480 ( .A1(n1843), .A2(n1321), .ZN(n987) );
  NAND2_X2 U2481 ( .A1(n998), .A2(n997), .ZN(n989) );
  NAND2_X2 U2482 ( .A1(n99), .A2(n988), .ZN(n992) );
  NOR2_X2 U2483 ( .A1(n995), .A2(n994), .ZN(n993) );
  NOR2_X2 U2484 ( .A1(n99), .A2(n3323), .ZN(n995) );
  XNOR2_X2 U2485 ( .A(n3468), .B(n3027), .ZN(n996) );
  NAND2_X2 U2486 ( .A1(n3311), .A2(n1217), .ZN(n997) );
  NAND2_X2 U2487 ( .A1(n58), .A2(n3310), .ZN(n998) );
  NAND2_X2 U2488 ( .A1(n999), .A2(n1602), .ZN(n1001) );
  INV_X2 U2489 ( .A(n1553), .ZN(n999) );
  INV_X2 U2490 ( .A(n2047), .ZN(n1325) );
  NAND2_X2 U2491 ( .A1(n1001), .A2(n1000), .ZN(n2047) );
  NAND2_X1 U2492 ( .A1(n1553), .A2(n2880), .ZN(n1000) );
  INV_X4 U2493 ( .A(n1002), .ZN(n2383) );
  NAND2_X2 U2494 ( .A1(n1006), .A2(n3095), .ZN(n1779) );
  NAND2_X2 U2498 ( .A1(n2383), .A2(n2087), .ZN(n1006) );
  NAND2_X2 U2499 ( .A1(n430), .A2(n1379), .ZN(n2087) );
  NOR2_X2 U2501 ( .A1(n1757), .A2(n1108), .ZN(n1002) );
  NAND2_X2 U2502 ( .A1(n681), .A2(n3106), .ZN(n1007) );
  NAND3_X2 U2503 ( .A1(n1744), .A2(n2232), .A3(n1795), .ZN(n1008) );
  NAND2_X2 U2504 ( .A1(n1010), .A2(n1009), .ZN(n2231) );
  INV_X2 U2506 ( .A(n3160), .ZN(n1012) );
  NOR2_X2 U2507 ( .A1(n2276), .A2(n2190), .ZN(n3162) );
  NAND2_X2 U2508 ( .A1(n1767), .A2(n3398), .ZN(n3420) );
  AOI22_X2 U2509 ( .A1(n1377), .A2(n2228), .B1(n4045), .B2(n93), .ZN(n2956) );
  BUF_X4 U2511 ( .A(n2332), .Z(n1016) );
  INV_X4 U2512 ( .A(n2332), .ZN(n3455) );
  NAND2_X2 U2514 ( .A1(n2050), .A2(n1019), .ZN(n1535) );
  NAND2_X2 U2515 ( .A1(n1171), .A2(n1170), .ZN(n2050) );
  AOI21_X2 U2518 ( .B1(n2395), .B2(n1022), .A(n1577), .ZN(n3102) );
  INV_X2 U2519 ( .A(n1022), .ZN(n3099) );
  NAND2_X1 U2520 ( .A1(n2167), .A2(n1022), .ZN(n1437) );
  NAND2_X2 U2521 ( .A1(n3404), .A2(n1025), .ZN(n2321) );
  NOR2_X2 U2523 ( .A1(n3040), .A2(n4178), .ZN(n1029) );
  INV_X2 U2525 ( .A(n1709), .ZN(n1030) );
  NAND2_X2 U2526 ( .A1(n1231), .A2(n1784), .ZN(n2897) );
  NOR2_X2 U2527 ( .A1(n2556), .A2(n3176), .ZN(n1766) );
  OAI21_X2 U2529 ( .B1(n3227), .B2(n4153), .A(n3228), .ZN(n1037) );
  INV_X4 U2530 ( .A(n3226), .ZN(n3227) );
  NAND2_X2 U2531 ( .A1(n1041), .A2(n1040), .ZN(n3576) );
  NAND2_X2 U2533 ( .A1(n1039), .A2(n2749), .ZN(n1041) );
  NAND2_X2 U2534 ( .A1(n2747), .A2(n2746), .ZN(n1039) );
  AOI22_X2 U2535 ( .A1(n2773), .A2(n2772), .B1(n2771), .B2(n2770), .ZN(n3377)
         );
  NAND3_X2 U2536 ( .A1(n2747), .A2(n2748), .A3(n2746), .ZN(n1040) );
  NAND2_X2 U2537 ( .A1(n2774), .A2(n2775), .ZN(n3375) );
  NAND2_X2 U2541 ( .A1(n1051), .A2(n1050), .ZN(n1811) );
  NAND2_X2 U2542 ( .A1(n2970), .A2(n2968), .ZN(n1050) );
  INV_X2 U2543 ( .A(n2968), .ZN(n1052) );
  INV_X2 U2544 ( .A(n1961), .ZN(n1054) );
  INV_X2 U2545 ( .A(n1811), .ZN(n1505) );
  NOR2_X2 U2546 ( .A1(n1056), .A2(n2801), .ZN(n1055) );
  NAND3_X2 U2548 ( .A1(n1818), .A2(n3129), .A3(n3118), .ZN(n2222) );
  NOR2_X2 U2549 ( .A1(n1060), .A2(n2295), .ZN(n1685) );
  NOR2_X2 U2550 ( .A1(n3314), .A2(n1062), .ZN(n1061) );
  NAND2_X2 U2551 ( .A1(n1064), .A2(n1063), .ZN(n1062) );
  NOR2_X2 U2552 ( .A1(n3044), .A2(n2345), .ZN(n1067) );
  NAND2_X2 U2553 ( .A1(n1659), .A2(n55), .ZN(n1891) );
  NAND2_X1 U2554 ( .A1(n1659), .A2(n3468), .ZN(n3410) );
  NAND2_X1 U2555 ( .A1(n1659), .A2(a[22]), .ZN(n1175) );
  NAND2_X2 U2556 ( .A1(n1353), .A2(n3183), .ZN(n3245) );
  INV_X4 U2557 ( .A(n1071), .ZN(n1616) );
  NOR2_X2 U2558 ( .A1(n1633), .A2(n3243), .ZN(n1071) );
  NAND2_X2 U2559 ( .A1(n1073), .A2(n1072), .ZN(n1633) );
  NOR2_X2 U2561 ( .A1(n1074), .A2(n827), .ZN(n2111) );
  NAND2_X2 U2562 ( .A1(n1074), .A2(n827), .ZN(n1124) );
  OAI21_X1 U2563 ( .B1(n4141), .B2(n1557), .A(n73), .ZN(n1075) );
  NAND3_X2 U2566 ( .A1(n1971), .A2(n1972), .A3(n1077), .ZN(n3434) );
  INV_X2 U2567 ( .A(n1078), .ZN(n1077) );
  NAND2_X2 U2568 ( .A1(n1080), .A2(n1079), .ZN(n1078) );
  NAND2_X1 U2569 ( .A1(n3455), .A2(n3534), .ZN(n1079) );
  NAND2_X1 U2570 ( .A1(n3454), .A2(a[3]), .ZN(n1080) );
  INV_X2 U2571 ( .A(n2120), .ZN(n3155) );
  NAND2_X2 U2572 ( .A1(n1083), .A2(n2120), .ZN(n3185) );
  NAND2_X2 U2573 ( .A1(n1082), .A2(n1081), .ZN(n2120) );
  XNOR2_X2 U2574 ( .A(n1913), .B(n2697), .ZN(n1082) );
  INV_X2 U2575 ( .A(n3148), .ZN(n1083) );
  NOR2_X2 U2576 ( .A1(n1084), .A2(n475), .ZN(n3148) );
  INV_X4 U2577 ( .A(n1360), .ZN(n1084) );
  NOR2_X2 U2578 ( .A1(n1953), .A2(n1947), .ZN(n1085) );
  INV_X2 U2579 ( .A(n1208), .ZN(n1947) );
  NAND2_X2 U2580 ( .A1(n1086), .A2(n1517), .ZN(n1953) );
  INV_X4 U2582 ( .A(n1087), .ZN(n2165) );
  BUF_X4 U2583 ( .A(n2384), .Z(n1088) );
  NAND3_X2 U2584 ( .A1(n1092), .A2(n1091), .A3(n1089), .ZN(n1456) );
  NAND2_X1 U2585 ( .A1(n1090), .A2(n2983), .ZN(n1089) );
  NOR2_X1 U2586 ( .A1(n91), .A2(n55), .ZN(n1090) );
  NAND2_X1 U2587 ( .A1(n2384), .A2(n2438), .ZN(n1091) );
  INV_X1 U2589 ( .A(n3334), .ZN(n1096) );
  NAND2_X2 U2590 ( .A1(n1093), .A2(n3334), .ZN(n1095) );
  NAND2_X2 U2591 ( .A1(n2364), .A2(n2363), .ZN(n1093) );
  NAND2_X2 U2592 ( .A1(n1095), .A2(n1094), .ZN(n3399) );
  INV_X2 U2593 ( .A(n3399), .ZN(n1097) );
  NAND2_X2 U2594 ( .A1(n2285), .A2(n2994), .ZN(n1574) );
  NAND2_X2 U2595 ( .A1(n1458), .A2(n1457), .ZN(n2994) );
  NOR3_X2 U2596 ( .A1(n1380), .A2(n1098), .A3(n2011), .ZN(n1540) );
  NAND2_X2 U2597 ( .A1(n1364), .A2(n1318), .ZN(n1098) );
  NAND2_X2 U2599 ( .A1(n3348), .A2(n3351), .ZN(n1101) );
  INV_X2 U2600 ( .A(n3297), .ZN(n3296) );
  INV_X2 U2601 ( .A(b[4]), .ZN(n2333) );
  NAND2_X2 U2602 ( .A1(n1104), .A2(n1103), .ZN(n1739) );
  NOR2_X2 U2603 ( .A1(n2169), .A2(n2171), .ZN(n1823) );
  NAND2_X2 U2604 ( .A1(n1107), .A2(n2216), .ZN(n2219) );
  NAND2_X2 U2605 ( .A1(n1734), .A2(n1733), .ZN(n1108) );
  NAND3_X2 U2606 ( .A1(n2293), .A2(n2097), .A3(n2904), .ZN(n1733) );
  NAND2_X2 U2608 ( .A1(n1110), .A2(n1109), .ZN(n1757) );
  NAND2_X2 U2609 ( .A1(n3085), .A2(n2046), .ZN(n1109) );
  AOI21_X2 U2611 ( .B1(n1454), .B2(n439), .A(n473), .ZN(n2116) );
  NAND2_X2 U2612 ( .A1(n1113), .A2(n2329), .ZN(n3567) );
  NOR2_X2 U2613 ( .A1(n1113), .A2(n2329), .ZN(n3564) );
  INV_X4 U2614 ( .A(n3298), .ZN(n1113) );
  NOR2_X2 U2619 ( .A1(n3109), .A2(n1121), .ZN(n2550) );
  NAND2_X2 U2622 ( .A1(n2868), .A2(n2869), .ZN(n1916) );
  NAND2_X2 U2625 ( .A1(n1625), .A2(n1624), .ZN(n1626) );
  NAND2_X2 U2626 ( .A1(n1127), .A2(n1126), .ZN(n1128) );
  NAND2_X1 U2627 ( .A1(n1382), .A2(n830), .ZN(n1126) );
  NAND2_X2 U2629 ( .A1(n1128), .A2(n1439), .ZN(n1532) );
  NAND2_X2 U2630 ( .A1(n3431), .A2(n3217), .ZN(n1130) );
  INV_X8 U2631 ( .A(n1131), .ZN(n2084) );
  NAND3_X2 U2632 ( .A1(n3633), .A2(n3632), .A3(n3634), .ZN(\d[33] ) );
  NAND2_X2 U2633 ( .A1(n3294), .A2(n1244), .ZN(n3295) );
  NAND2_X2 U2634 ( .A1(n1451), .A2(n1450), .ZN(n1244) );
  NAND2_X4 U2635 ( .A1(n1514), .A2(n1513), .ZN(n3294) );
  NAND2_X2 U2636 ( .A1(n3249), .A2(n3293), .ZN(n2003) );
  NAND2_X2 U2638 ( .A1(n1137), .A2(n1997), .ZN(n2583) );
  INV_X2 U2639 ( .A(n2464), .ZN(n1137) );
  NAND2_X2 U2642 ( .A1(n1140), .A2(n2476), .ZN(n1405) );
  INV_X1 U2645 ( .A(n1143), .ZN(n1142) );
  AOI21_X1 U2646 ( .B1(n1144), .B2(n3529), .A(n3507), .ZN(n1143) );
  INV_X1 U2647 ( .A(n1154), .ZN(n1144) );
  NAND2_X1 U2648 ( .A1(n1148), .A2(n1146), .ZN(n1145) );
  NAND3_X1 U2649 ( .A1(n1147), .A2(n1153), .A3(n1154), .ZN(n1146) );
  INV_X1 U2650 ( .A(n3529), .ZN(n1147) );
  INV_X1 U2651 ( .A(n1153), .ZN(n1149) );
  OAI22_X1 U2652 ( .A1(n3527), .A2(n455), .B1(n3532), .B2(n3500), .ZN(n1153)
         );
  AOI21_X2 U2653 ( .B1(n1784), .B2(n1235), .A(n1150), .ZN(n3529) );
  AOI22_X1 U2656 ( .A1(n3497), .A2(n3500), .B1(n3532), .B2(n3528), .ZN(n1154)
         );
  NAND2_X2 U2657 ( .A1(b[11]), .A2(b[12]), .ZN(n3009) );
  INV_X2 U2659 ( .A(n2605), .ZN(n1155) );
  NAND2_X2 U2660 ( .A1(n2604), .A2(n2605), .ZN(n1156) );
  NAND2_X2 U2661 ( .A1(n1158), .A2(n1157), .ZN(n2504) );
  INV_X2 U2662 ( .A(n1159), .ZN(n1158) );
  NAND2_X2 U2664 ( .A1(n1873), .A2(n2504), .ZN(n2492) );
  NAND2_X2 U2665 ( .A1(n2485), .A2(n2484), .ZN(n1873) );
  NOR2_X1 U2666 ( .A1(n3083), .A2(n1160), .ZN(n3356) );
  NAND2_X1 U2667 ( .A1(n3083), .A2(n1160), .ZN(n3357) );
  INV_X2 U2668 ( .A(n1576), .ZN(n3777) );
  NAND2_X2 U2669 ( .A1(n2173), .A2(n2172), .ZN(n1576) );
  NAND2_X2 U2670 ( .A1(n1271), .A2(n3777), .ZN(n3556) );
  NAND2_X2 U2671 ( .A1(n1803), .A2(n964), .ZN(n1271) );
  NAND3_X2 U2672 ( .A1(n1289), .A2(n3383), .A3(n3382), .ZN(n2172) );
  NAND2_X2 U2673 ( .A1(n1161), .A2(n2943), .ZN(n3171) );
  INV_X4 U2674 ( .A(b[7]), .ZN(n1597) );
  INV_X4 U2677 ( .A(n1163), .ZN(n2931) );
  NOR2_X4 U2678 ( .A1(n1164), .A2(n2777), .ZN(n1292) );
  AOI21_X2 U2679 ( .B1(n1359), .B2(n1358), .A(n91), .ZN(n1164) );
  NAND2_X1 U2682 ( .A1(n1750), .A2(n1168), .ZN(n1746) );
  NOR2_X1 U2683 ( .A1(n1750), .A2(n1168), .ZN(n1747) );
  XNOR2_X2 U2684 ( .A(n1750), .B(n1168), .ZN(n1749) );
  AOI21_X2 U2685 ( .B1(n3430), .B2(n2998), .A(n4085), .ZN(n1168) );
  INV_X1 U2686 ( .A(n2207), .ZN(n2565) );
  NAND3_X2 U2687 ( .A1(n3733), .A2(n3731), .A3(n3732), .ZN(\d[34] ) );
  INV_X4 U2688 ( .A(n1832), .ZN(n2386) );
  BUF_X4 U2693 ( .A(n1687), .Z(n1180) );
  INV_X2 U2695 ( .A(n2967), .ZN(n2971) );
  NAND2_X2 U2697 ( .A1(n1187), .A2(n2593), .ZN(n1188) );
  NAND2_X2 U2698 ( .A1(n2589), .A2(n2394), .ZN(n1187) );
  NAND2_X2 U2699 ( .A1(n4072), .A2(n3982), .ZN(\d[20]_BAR ) );
  NAND3_X2 U2701 ( .A1(n1196), .A2(n1194), .A3(n1193), .ZN(n3064) );
  NAND3_X2 U2702 ( .A1(n3056), .A2(n1195), .A3(n3055), .ZN(n1194) );
  INV_X1 U2703 ( .A(n3054), .ZN(n1195) );
  INV_X2 U2705 ( .A(n2929), .ZN(n2926) );
  NAND3_X2 U2706 ( .A1(n2838), .A2(n2837), .A3(n2387), .ZN(n2839) );
  NAND2_X2 U2707 ( .A1(n2835), .A2(n2834), .ZN(n2840) );
  INV_X1 U2708 ( .A(n2905), .ZN(n2097) );
  OAI21_X2 U2709 ( .B1(n2874), .B2(n2881), .A(n2873), .ZN(n2905) );
  NAND2_X2 U2710 ( .A1(n1199), .A2(n3357), .ZN(n3359) );
  INV_X2 U2711 ( .A(n3356), .ZN(n1199) );
  NOR2_X2 U2712 ( .A1(n3082), .A2(n3081), .ZN(n3083) );
  INV_X2 U2713 ( .A(n3257), .ZN(n3256) );
  NAND2_X2 U2714 ( .A1(n1201), .A2(n1200), .ZN(n2190) );
  NOR2_X2 U2717 ( .A1(n2914), .A2(n2177), .ZN(n2945) );
  NOR2_X1 U2718 ( .A1(n3814), .A2(n3798), .ZN(n3789) );
  INV_X1 U2722 ( .A(n3582), .ZN(n3585) );
  NAND2_X2 U2723 ( .A1(n2384), .A2(n54), .ZN(n2298) );
  NAND2_X2 U2724 ( .A1(n2856), .A2(n2855), .ZN(n1812) );
  INV_X4 U2725 ( .A(n2069), .ZN(n3266) );
  AOI21_X1 U2726 ( .B1(n86), .B2(a[8]), .A(n1993), .ZN(n1992) );
  NAND2_X1 U2727 ( .A1(n86), .A2(n93), .ZN(n2243) );
  OAI21_X1 U2731 ( .B1(n3262), .B2(n3261), .A(n3260), .ZN(n3281) );
  NAND2_X2 U2733 ( .A1(n2294), .A2(n3266), .ZN(n1226) );
  NOR2_X4 U2734 ( .A1(n2664), .A2(n2663), .ZN(n2760) );
  NAND2_X2 U2735 ( .A1(n2383), .A2(n2087), .ZN(n1207) );
  NOR2_X2 U2737 ( .A1(n2503), .A2(n2490), .ZN(n2491) );
  INV_X8 U2738 ( .A(n3460), .ZN(n1209) );
  NAND2_X1 U2739 ( .A1(n10), .A2(n64), .ZN(n3175) );
  NAND2_X2 U2742 ( .A1(n3328), .A2(n100), .ZN(n1215) );
  NAND2_X1 U2743 ( .A1(n2084), .A2(n3468), .ZN(n1216) );
  NAND2_X2 U2744 ( .A1(n1215), .A2(n1216), .ZN(n2887) );
  BUF_X4 U2745 ( .A(n3475), .Z(n1217) );
  NAND2_X1 U2747 ( .A1(n1287), .A2(n4064), .ZN(n1219) );
  INV_X4 U2748 ( .A(n58), .ZN(n1221) );
  NOR2_X2 U2749 ( .A1(n2979), .A2(n2978), .ZN(n2993) );
  NAND2_X2 U2750 ( .A1(n3573), .A2(n3574), .ZN(n1850) );
  AOI22_X2 U2751 ( .A1(n3010), .A2(n3178), .B1(n1837), .B2(n3179), .ZN(n1880)
         );
  NAND2_X1 U2752 ( .A1(n3177), .A2(n2228), .ZN(n3178) );
  NOR2_X4 U2753 ( .A1(n2083), .A2(n3154), .ZN(n2082) );
  INV_X1 U2755 ( .A(n1602), .ZN(n1224) );
  NAND2_X2 U2757 ( .A1(n2711), .A2(n2710), .ZN(n2713) );
  NAND2_X2 U2758 ( .A1(n1893), .A2(n743), .ZN(n1356) );
  NAND2_X2 U2759 ( .A1(n1654), .A2(n1653), .ZN(n1230) );
  NAND2_X2 U2760 ( .A1(n1654), .A2(n1653), .ZN(n2962) );
  INV_X1 U2761 ( .A(n1449), .ZN(n3430) );
  NAND2_X2 U2762 ( .A1(n2091), .A2(n1495), .ZN(n2090) );
  NOR2_X2 U2763 ( .A1(n3192), .A2(n21), .ZN(n2080) );
  INV_X2 U2764 ( .A(n2433), .ZN(n1567) );
  NOR2_X1 U2766 ( .A1(n3659), .A2(n3658), .ZN(n3663) );
  NOR3_X1 U2767 ( .A1(n3615), .A2(n3675), .A3(n3659), .ZN(n3616) );
  INV_X2 U2768 ( .A(n70), .ZN(n1233) );
  INV_X1 U2769 ( .A(n2368), .ZN(n1234) );
  NAND3_X2 U2770 ( .A1(n2235), .A2(n2278), .A3(n3193), .ZN(n2233) );
  INV_X2 U2771 ( .A(n1407), .ZN(n1235) );
  NOR2_X4 U2772 ( .A1(n3241), .A2(n2063), .ZN(n3242) );
  NOR2_X4 U2773 ( .A1(n3736), .A2(n3737), .ZN(n3947) );
  INV_X4 U2774 ( .A(n2354), .ZN(n1237) );
  NOR2_X2 U2775 ( .A1(n3136), .A2(n3137), .ZN(n1238) );
  INV_X1 U2776 ( .A(n1238), .ZN(n3152) );
  INV_X2 U2777 ( .A(n3184), .ZN(n1343) );
  INV_X2 U2779 ( .A(n3229), .ZN(n3232) );
  NAND2_X2 U2781 ( .A1(n1239), .A2(n1240), .ZN(n1242) );
  INV_X2 U2782 ( .A(n3353), .ZN(n1239) );
  NAND2_X2 U2784 ( .A1(n2299), .A2(n2300), .ZN(n2161) );
  INV_X1 U2785 ( .A(n3059), .ZN(n3060) );
  NAND2_X2 U2786 ( .A1(n1616), .A2(n1615), .ZN(n2103) );
  NAND2_X2 U2787 ( .A1(n3794), .A2(n466), .ZN(n1243) );
  NAND2_X2 U2788 ( .A1(n3151), .A2(n3150), .ZN(n3157) );
  NAND2_X1 U2791 ( .A1(n2045), .A2(n2299), .ZN(n3517) );
  NAND2_X2 U2794 ( .A1(n3318), .A2(n3317), .ZN(n3348) );
  NAND2_X1 U2796 ( .A1(n2157), .A2(n1784), .ZN(n2156) );
  NAND2_X1 U2797 ( .A1(n2758), .A2(n2757), .ZN(n1250) );
  NAND2_X2 U2799 ( .A1(n1250), .A2(n1251), .ZN(n2665) );
  NAND2_X1 U2803 ( .A1(n2665), .A2(n2760), .ZN(n1255) );
  NAND2_X2 U2804 ( .A1(n1255), .A2(n1256), .ZN(n1452) );
  INV_X1 U2805 ( .A(n2665), .ZN(n1254) );
  INV_X1 U2806 ( .A(n1319), .ZN(n1257) );
  NAND2_X2 U2807 ( .A1(n3216), .A2(n3215), .ZN(n3259) );
  NOR3_X2 U2808 ( .A1(n3870), .A2(n3871), .A3(n3872), .ZN(n3881) );
  NOR2_X2 U2809 ( .A1(n1509), .A2(n2237), .ZN(n2236) );
  BUF_X4 U2810 ( .A(n3455), .Z(n1262) );
  NOR2_X2 U2813 ( .A1(n22), .A2(n4008), .ZN(n1618) );
  NAND2_X1 U2814 ( .A1(n2584), .A2(n2647), .ZN(n1268) );
  NAND2_X2 U2816 ( .A1(n1561), .A2(n1562), .ZN(n1272) );
  NAND3_X2 U2817 ( .A1(n3557), .A2(n2012), .A3(n1408), .ZN(n1273) );
  NAND2_X1 U2818 ( .A1(n3718), .A2(n3716), .ZN(n3717) );
  NAND2_X2 U2819 ( .A1(n1274), .A2(n1275), .ZN(n3087) );
  NAND2_X2 U2821 ( .A1(n1277), .A2(n81), .ZN(n1279) );
  NOR2_X2 U2822 ( .A1(n1480), .A2(n2869), .ZN(n1280) );
  NAND2_X2 U2824 ( .A1(n2229), .A2(n3057), .ZN(n1726) );
  NAND2_X2 U2825 ( .A1(n1209), .A2(a[10]), .ZN(n2229) );
  NAND2_X2 U2828 ( .A1(n3180), .A2(n3185), .ZN(n3246) );
  NAND2_X1 U2829 ( .A1(n3830), .A2(n3904), .ZN(n3832) );
  NAND2_X4 U2830 ( .A1(n2118), .A2(n2067), .ZN(n4003) );
  INV_X4 U2831 ( .A(n4018), .ZN(n1482) );
  NAND2_X1 U2833 ( .A1(n3292), .A2(n3291), .ZN(n1283) );
  NOR2_X2 U2834 ( .A1(n3963), .A2(n22), .ZN(n3970) );
  NOR2_X2 U2835 ( .A1(n3542), .A2(n1665), .ZN(n1664) );
  INV_X1 U2836 ( .A(n1678), .ZN(n1665) );
  NOR2_X1 U2837 ( .A1(n3192), .A2(n21), .ZN(n1285) );
  INV_X4 U2838 ( .A(n3205), .ZN(n1301) );
  NAND2_X2 U2839 ( .A1(n4166), .A2(n1611), .ZN(n1287) );
  NAND2_X2 U2840 ( .A1(n3431), .A2(n3109), .ZN(n3111) );
  NAND2_X2 U2841 ( .A1(n2236), .A2(n1601), .ZN(n1288) );
  NAND2_X2 U2842 ( .A1(n1601), .A2(n2236), .ZN(n3605) );
  NAND2_X2 U2843 ( .A1(n3322), .A2(n3321), .ZN(n1289) );
  OAI21_X2 U2844 ( .B1(n3058), .B2(n3054), .A(n3012), .ZN(n1290) );
  INV_X1 U2846 ( .A(n2512), .ZN(n1291) );
  INV_X2 U2847 ( .A(n3558), .ZN(n3788) );
  NAND2_X1 U2848 ( .A1(n3311), .A2(n97), .ZN(n1825) );
  NAND2_X1 U2850 ( .A1(n3402), .A2(n3403), .ZN(n1692) );
  INV_X4 U2851 ( .A(n3427), .ZN(n3311) );
  NOR2_X1 U2852 ( .A1(n1370), .A2(n3534), .ZN(n2292) );
  NOR2_X1 U2853 ( .A1(n1370), .A2(n3407), .ZN(n2322) );
  NOR3_X2 U2854 ( .A1(n3536), .A2(n2292), .A3(n2291), .ZN(n3550) );
  NAND2_X2 U2855 ( .A1(n2042), .A2(n2041), .ZN(n2104) );
  NAND2_X2 U2857 ( .A1(n1600), .A2(b[11]), .ZN(n3205) );
  NAND2_X1 U2858 ( .A1(n1790), .A2(n2768), .ZN(n1296) );
  INV_X2 U2860 ( .A(n1790), .ZN(n1294) );
  INV_X1 U2861 ( .A(n2768), .ZN(n1295) );
  INV_X4 U2863 ( .A(n3085), .ZN(n1417) );
  AOI21_X1 U2864 ( .B1(n2992), .B2(n2976), .A(n2975), .ZN(n1507) );
  INV_X4 U2866 ( .A(n2282), .ZN(n2281) );
  NOR2_X4 U2867 ( .A1(n2987), .A2(n2986), .ZN(n2282) );
  AOI22_X2 U2869 ( .A1(n3053), .A2(n1728), .B1(n83), .B2(n3052), .ZN(n1298) );
  INV_X8 U2871 ( .A(n1301), .ZN(n1303) );
  INV_X2 U2872 ( .A(n1223), .ZN(n1853) );
  NAND2_X2 U2873 ( .A1(n1432), .A2(n1433), .ZN(n1435) );
  NAND3_X2 U2874 ( .A1(n2034), .A2(n2033), .A3(n2032), .ZN(n1304) );
  OAI21_X1 U2875 ( .B1(n3398), .B2(n3400), .A(n3399), .ZN(n3336) );
  NAND2_X2 U2879 ( .A1(n3990), .A2(n3933), .ZN(n1309) );
  NAND2_X2 U2880 ( .A1(n3990), .A2(n3933), .ZN(n3994) );
  OAI21_X1 U2881 ( .B1(n1314), .B2(n3362), .A(n3361), .ZN(n1310) );
  INV_X1 U2882 ( .A(n3058), .ZN(n3056) );
  NAND2_X2 U2883 ( .A1(n1912), .A2(n4150), .ZN(n1529) );
  NAND2_X2 U2884 ( .A1(n1984), .A2(n1989), .ZN(n1311) );
  INV_X1 U2886 ( .A(n3814), .ZN(n1312) );
  NAND2_X2 U2887 ( .A1(n4155), .A2(n3007), .ZN(n1313) );
  NAND2_X2 U2888 ( .A1(n4155), .A2(n3007), .ZN(n3013) );
  INV_X4 U2889 ( .A(n2286), .ZN(n1319) );
  NOR2_X2 U2890 ( .A1(n1464), .A2(n1844), .ZN(n1314) );
  INV_X4 U2891 ( .A(n3981), .ZN(n1320) );
  NAND2_X1 U2892 ( .A1(n1784), .A2(n3453), .ZN(n1972) );
  NAND2_X2 U2893 ( .A1(b[8]), .A2(b[7]), .ZN(n1598) );
  NAND2_X2 U2894 ( .A1(n2962), .A2(n18), .ZN(n2277) );
  NAND2_X4 U2895 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
  INV_X1 U2896 ( .A(n2014), .ZN(n1322) );
  AOI22_X2 U2897 ( .A1(n3153), .A2(n3157), .B1(n3180), .B2(n3155), .ZN(n2083)
         );
  INV_X4 U2898 ( .A(b[9]), .ZN(n1323) );
  INV_X4 U2899 ( .A(b[9]), .ZN(n2423) );
  NAND2_X1 U2900 ( .A1(n3120), .A2(n88), .ZN(n1327) );
  INV_X4 U2904 ( .A(n2912), .ZN(n2911) );
  NAND2_X2 U2905 ( .A1(n2910), .A2(n2911), .ZN(n1684) );
  NAND2_X2 U2906 ( .A1(n2058), .A2(n37), .ZN(n1330) );
  AOI21_X2 U2907 ( .B1(n2651), .B2(n2650), .A(n2649), .ZN(n2676) );
  INV_X4 U2908 ( .A(n3419), .ZN(n1551) );
  NAND2_X1 U2909 ( .A1(n99), .A2(n3431), .ZN(n1660) );
  AOI22_X2 U2911 ( .A1(n1988), .A2(n1987), .B1(n1986), .B2(n1985), .ZN(n3608)
         );
  NAND2_X2 U2912 ( .A1(n4003), .A2(n4004), .ZN(n1623) );
  NAND2_X2 U2913 ( .A1(n2511), .A2(n2510), .ZN(n1334) );
  NAND2_X2 U2914 ( .A1(n1332), .A2(n1333), .ZN(n1335) );
  XNOR2_X2 U2917 ( .A(n3287), .B(n69), .ZN(n1939) );
  INV_X4 U2920 ( .A(n1227), .ZN(n2299) );
  NAND2_X1 U2922 ( .A1(n3184), .A2(n3159), .ZN(n1344) );
  OAI21_X1 U2925 ( .B1(n3622), .B2(n3667), .A(n3621), .ZN(n3623) );
  INV_X1 U2926 ( .A(n3667), .ZN(n3670) );
  AOI21_X2 U2927 ( .B1(n1998), .B2(n2598), .A(n2597), .ZN(n2626) );
  NAND2_X2 U2928 ( .A1(n1612), .A2(n1611), .ZN(n2930) );
  NAND3_X1 U2929 ( .A1(n4047), .A2(n1996), .A3(n1994), .ZN(n1346) );
  NAND2_X2 U2931 ( .A1(n2368), .A2(n70), .ZN(n1446) );
  NAND2_X2 U2932 ( .A1(n666), .A2(n1965), .ZN(n1350) );
  INV_X2 U2933 ( .A(n1969), .ZN(n1351) );
  INV_X1 U2934 ( .A(n3451), .ZN(n1352) );
  INV_X1 U2935 ( .A(n2445), .ZN(n2340) );
  NAND2_X2 U2936 ( .A1(n2445), .A2(n2302), .ZN(n2514) );
  XNOR2_X1 U2937 ( .A(n2320), .B(n3805), .ZN(n3807) );
  XNOR2_X2 U2938 ( .A(n2585), .B(n2588), .ZN(n2499) );
  NAND2_X1 U2939 ( .A1(n4045), .A2(a[19]), .ZN(n2450) );
  NAND2_X2 U2940 ( .A1(n3745), .A2(n3813), .ZN(n2269) );
  INV_X4 U2941 ( .A(n2527), .ZN(n1893) );
  NAND2_X2 U2942 ( .A1(n1357), .A2(n98), .ZN(n1359) );
  INV_X2 U2943 ( .A(n1913), .ZN(n1357) );
  NOR2_X4 U2944 ( .A1(n2122), .A2(n1942), .ZN(n2063) );
  NOR2_X1 U2945 ( .A1(n3954), .A2(n4008), .ZN(n3971) );
  NOR2_X1 U2946 ( .A1(n43), .A2(n3762), .ZN(n3764) );
  AOI21_X1 U2947 ( .B1(n43), .B2(n3762), .A(n3761), .ZN(n3765) );
  INV_X1 U2948 ( .A(n3734), .ZN(n3604) );
  NOR3_X1 U2949 ( .A1(n3852), .A2(n854), .A3(n3853), .ZN(n3861) );
  INV_X2 U2950 ( .A(n3252), .ZN(n1366) );
  INV_X2 U2951 ( .A(n2321), .ZN(n1369) );
  INV_X4 U2953 ( .A(n1271), .ZN(n1829) );
  INV_X4 U2954 ( .A(n2082), .ZN(n2033) );
  NOR2_X2 U2955 ( .A1(n3158), .A2(n3191), .ZN(n2032) );
  INV_X1 U2956 ( .A(n2952), .ZN(n2951) );
  INV_X1 U2957 ( .A(n3203), .ZN(n2157) );
  NAND2_X1 U2958 ( .A1(n249), .A2(n56), .ZN(n3141) );
  NAND2_X1 U2960 ( .A1(n2530), .A2(n2531), .ZN(n2532) );
  NAND2_X2 U2961 ( .A1(n2529), .A2(n1991), .ZN(n1499) );
  INV_X8 U2962 ( .A(n3080), .ZN(n1377) );
  NAND2_X4 U2963 ( .A1(n1613), .A2(n1614), .ZN(n2125) );
  NAND2_X1 U2964 ( .A1(n2563), .A2(n2562), .ZN(n3273) );
  NAND2_X2 U2965 ( .A1(n1502), .A2(n1590), .ZN(n1380) );
  BUF_X4 U2966 ( .A(n2084), .Z(n1381) );
  INV_X1 U2968 ( .A(n2917), .ZN(n2915) );
  NOR2_X2 U2969 ( .A1(n2242), .A2(n441), .ZN(n2917) );
  XNOR2_X2 U2970 ( .A(n3251), .B(n3250), .ZN(n3252) );
  NAND2_X2 U2971 ( .A1(n3076), .A2(n3075), .ZN(n3077) );
  NAND2_X1 U2974 ( .A1(n1617), .A2(n3970), .ZN(n3965) );
  INV_X1 U2975 ( .A(n2953), .ZN(n2955) );
  INV_X1 U2976 ( .A(n3305), .ZN(n2367) );
  NAND2_X1 U2977 ( .A1(n1980), .A2(n3275), .ZN(n1385) );
  NAND2_X2 U2978 ( .A1(n1209), .A2(n3124), .ZN(n2175) );
  NAND2_X1 U2979 ( .A1(n2980), .A2(n54), .ZN(n1387) );
  NAND2_X1 U2980 ( .A1(n2022), .A2(n97), .ZN(n1388) );
  NAND2_X1 U2981 ( .A1(n1387), .A2(n1388), .ZN(n2578) );
  INV_X4 U2982 ( .A(n1833), .ZN(n1559) );
  NAND2_X2 U2983 ( .A1(n2386), .A2(n2891), .ZN(n1390) );
  NOR2_X2 U2985 ( .A1(n2080), .A2(n3191), .ZN(n2038) );
  INV_X4 U2987 ( .A(n3106), .ZN(n1744) );
  INV_X1 U2990 ( .A(n3550), .ZN(n3551) );
  NOR2_X1 U2991 ( .A1(n4167), .A2(n3550), .ZN(n3553) );
  INV_X1 U2994 ( .A(n1396), .ZN(n3471) );
  XOR2_X2 U2995 ( .A(n3465), .B(n3466), .Z(n1397) );
  INV_X4 U2996 ( .A(n2039), .ZN(n1877) );
  NAND2_X1 U2997 ( .A1(n3718), .A2(n3721), .ZN(n3725) );
  NAND2_X2 U2998 ( .A1(n1581), .A2(n1582), .ZN(n1400) );
  NAND2_X4 U3000 ( .A1(n3572), .A2(n1639), .ZN(n1938) );
  OAI21_X1 U3001 ( .B1(n3719), .B2(n3718), .A(n3717), .ZN(n3724) );
  INV_X1 U3002 ( .A(n2568), .ZN(n1404) );
  NAND3_X1 U3004 ( .A1(n3848), .A2(n3857), .A3(n4021), .ZN(n3862) );
  NAND2_X4 U3006 ( .A1(n2199), .A2(n2200), .ZN(n1449) );
  INV_X4 U3007 ( .A(n2238), .ZN(n1408) );
  NAND2_X1 U3010 ( .A1(n3379), .A2(n3378), .ZN(n1412) );
  INV_X2 U3011 ( .A(n3379), .ZN(n1411) );
  NAND2_X1 U3013 ( .A1(n3399), .A2(n3398), .ZN(n1415) );
  NAND2_X2 U3015 ( .A1(n1833), .A2(n3400), .ZN(n1561) );
  INV_X4 U3017 ( .A(n2046), .ZN(n1416) );
  NOR2_X1 U3019 ( .A1(n22), .A2(n1510), .ZN(n3742) );
  NAND2_X1 U3020 ( .A1(n2053), .A2(n3053), .ZN(n1423) );
  NAND2_X2 U3021 ( .A1(n1421), .A2(n1422), .ZN(n1424) );
  INV_X2 U3022 ( .A(n2053), .ZN(n1421) );
  NAND2_X2 U3024 ( .A1(n83), .A2(n1729), .ZN(n1426) );
  NAND2_X2 U3025 ( .A1(n1425), .A2(n1426), .ZN(n2053) );
  INV_X1 U3026 ( .A(n3362), .ZN(n1427) );
  OAI21_X2 U3027 ( .B1(n3329), .B2(n3538), .A(n3328), .ZN(n3403) );
  INV_X1 U3029 ( .A(n3185), .ZN(n3187) );
  NAND2_X2 U3030 ( .A1(n68), .A2(n3094), .ZN(n1429) );
  NAND2_X1 U3032 ( .A1(n3403), .A2(n3401), .ZN(n3330) );
  NAND2_X1 U3033 ( .A1(n2630), .A2(n1348), .ZN(n1434) );
  NAND2_X2 U3035 ( .A1(n1436), .A2(n3099), .ZN(n1438) );
  INV_X1 U3036 ( .A(n1531), .ZN(n1439) );
  NOR2_X1 U3037 ( .A1(n1309), .A2(n3993), .ZN(n3998) );
  AOI21_X2 U3038 ( .B1(n260), .B2(n2280), .A(n2279), .ZN(n2067) );
  NAND2_X1 U3039 ( .A1(n3939), .A2(n3940), .ZN(n3941) );
  NOR2_X1 U3040 ( .A1(n3907), .A2(n3906), .ZN(n3908) );
  NAND2_X2 U3042 ( .A1(n1443), .A2(n1442), .ZN(n1696) );
  XOR2_X1 U3043 ( .A(n3498), .B(a[24]), .Z(n2440) );
  NAND3_X1 U3044 ( .A1(n3066), .A2(n3498), .A3(n3413), .ZN(n3069) );
  NAND3_X1 U3045 ( .A1(n2333), .A2(n2145), .A3(n3498), .ZN(n2806) );
  INV_X2 U3046 ( .A(n3387), .ZN(n1444) );
  INV_X2 U3047 ( .A(n1745), .ZN(n1447) );
  INV_X2 U3048 ( .A(n3920), .ZN(n3873) );
  NAND3_X2 U3049 ( .A1(n2412), .A2(n2316), .A3(n1315), .ZN(n1448) );
  INV_X4 U3052 ( .A(n1452), .ZN(n2771) );
  NOR2_X2 U3053 ( .A1(n1418), .A2(n3823), .ZN(n3906) );
  NAND3_X1 U3054 ( .A1(n1088), .A2(n2045), .A3(n1645), .ZN(n3516) );
  INV_X1 U3055 ( .A(n1645), .ZN(n1453) );
  NOR2_X2 U3056 ( .A1(n86), .A2(n3139), .ZN(n2821) );
  OAI21_X1 U3057 ( .B1(n3078), .B2(n3079), .A(n3300), .ZN(n3358) );
  NAND2_X2 U3058 ( .A1(n1287), .A2(n4064), .ZN(n2137) );
  AOI21_X2 U3059 ( .B1(n2101), .B2(n3034), .A(n1880), .ZN(n3237) );
  NAND2_X2 U3060 ( .A1(n2198), .A2(a[17]), .ZN(n1555) );
  NAND2_X2 U3061 ( .A1(n2567), .A2(n2568), .ZN(n2310) );
  NAND2_X1 U3062 ( .A1(n2407), .A2(n2359), .ZN(n2318) );
  NAND2_X1 U3063 ( .A1(n1463), .A2(n2757), .ZN(n1462) );
  NAND2_X2 U3064 ( .A1(n2658), .A2(n2657), .ZN(n1463) );
  NAND2_X2 U3065 ( .A1(n3064), .A2(n3063), .ZN(n1464) );
  INV_X2 U3066 ( .A(n2186), .ZN(n1465) );
  INV_X4 U3067 ( .A(n2595), .ZN(n1998) );
  NAND2_X1 U3068 ( .A1(n1874), .A2(n201), .ZN(n1469) );
  NAND2_X2 U3069 ( .A1(n1469), .A2(n1470), .ZN(n3085) );
  NAND2_X2 U3071 ( .A1(n3243), .A2(n1633), .ZN(n1615) );
  INV_X4 U3073 ( .A(n2625), .ZN(n1943) );
  INV_X4 U3075 ( .A(n3236), .ZN(n1745) );
  NOR2_X2 U3076 ( .A1(n1273), .A2(n1260), .ZN(n1471) );
  NAND2_X2 U3077 ( .A1(n1472), .A2(n1473), .ZN(n3346) );
  NOR2_X2 U3079 ( .A1(n3420), .A2(n1552), .ZN(n3396) );
  NAND2_X4 U3080 ( .A1(n2000), .A2(n1999), .ZN(n2247) );
  NAND2_X2 U3082 ( .A1(n2151), .A2(n4068), .ZN(n1475) );
  INV_X4 U3083 ( .A(n1292), .ZN(n2139) );
  INV_X2 U3085 ( .A(n2844), .ZN(n1476) );
  INV_X1 U3086 ( .A(n2928), .ZN(n1477) );
  INV_X4 U3087 ( .A(n2556), .ZN(n1478) );
  OAI21_X1 U3089 ( .B1(n3929), .B2(n3602), .A(n3601), .ZN(n3625) );
  INV_X4 U3090 ( .A(n3129), .ZN(n3132) );
  INV_X4 U3091 ( .A(n3132), .ZN(n1487) );
  NAND2_X1 U3092 ( .A1(n1350), .A2(n1657), .ZN(n3779) );
  NAND2_X1 U3094 ( .A1(n3471), .A2(n3479), .ZN(n3480) );
  NAND2_X2 U3095 ( .A1(n2697), .A2(n3200), .ZN(n2204) );
  INV_X1 U3096 ( .A(n3806), .ZN(n1802) );
  AOI21_X1 U3097 ( .B1(n3358), .B2(n3357), .A(n3356), .ZN(n3362) );
  NAND2_X2 U3098 ( .A1(n2955), .A2(n2954), .ZN(n3164) );
  NAND2_X1 U3099 ( .A1(n3204), .A2(n3468), .ZN(n2793) );
  NAND2_X2 U3100 ( .A1(n1580), .A2(n2148), .ZN(n1581) );
  INV_X1 U3101 ( .A(n3022), .ZN(n1934) );
  INV_X4 U3103 ( .A(b[1]), .ZN(n2174) );
  NAND2_X1 U3104 ( .A1(n2404), .A2(n733), .ZN(n1484) );
  NAND2_X2 U3105 ( .A1(n1484), .A2(n1485), .ZN(n2102) );
  NAND2_X1 U3106 ( .A1(n95), .A2(n3200), .ZN(n1975) );
  OR2_X4 U3107 ( .A1(n2155), .A2(n1236), .ZN(n1486) );
  NOR2_X1 U3110 ( .A1(n3303), .A2(a[7]), .ZN(n3414) );
  NOR2_X1 U3111 ( .A1(n3186), .A2(n3152), .ZN(n3153) );
  NAND2_X1 U3112 ( .A1(n2579), .A2(n53), .ZN(n1490) );
  INV_X4 U3113 ( .A(n2785), .ZN(n2334) );
  NOR2_X4 U3114 ( .A1(n1568), .A2(n2125), .ZN(n2069) );
  NAND2_X2 U3115 ( .A1(n2925), .A2(n1292), .ZN(n1611) );
  NOR2_X1 U3116 ( .A1(n3788), .A2(n3787), .ZN(n3798) );
  NAND2_X2 U3117 ( .A1(n2447), .A2(n2448), .ZN(n2501) );
  NOR3_X1 U3118 ( .A1(n3714), .A2(n3660), .A3(n3709), .ZN(n3848) );
  INV_X1 U3119 ( .A(n3714), .ZN(n3715) );
  INV_X1 U3120 ( .A(n2672), .ZN(n2673) );
  INV_X1 U3121 ( .A(n2632), .ZN(n2635) );
  NAND2_X1 U3123 ( .A1(n1361), .A2(n2258), .ZN(n1493) );
  NAND2_X1 U3124 ( .A1(n3203), .A2(a[11]), .ZN(n1494) );
  INV_X2 U3125 ( .A(n62), .ZN(n1495) );
  NAND2_X2 U3126 ( .A1(n2492), .A2(n2491), .ZN(n1496) );
  NAND2_X2 U3127 ( .A1(n1318), .A2(n1364), .ZN(n1497) );
  NAND2_X2 U3128 ( .A1(n1499), .A2(n1500), .ZN(n2533) );
  INV_X4 U3129 ( .A(n2206), .ZN(n2205) );
  BUF_X4 U3131 ( .A(a[5]), .Z(n3475) );
  INV_X2 U3132 ( .A(n3352), .ZN(n3355) );
  NAND2_X2 U3134 ( .A1(n1579), .A2(n1384), .ZN(n1582) );
  NAND2_X1 U3135 ( .A1(n2195), .A2(n3560), .ZN(n2194) );
  NOR3_X1 U3137 ( .A1(n3067), .A2(n2506), .A3(a[12]), .ZN(n2883) );
  XNOR2_X1 U3142 ( .A(n2506), .B(a[25]), .ZN(n2476) );
  NAND2_X1 U3143 ( .A1(n1811), .A2(n2967), .ZN(n1506) );
  NOR2_X2 U3144 ( .A1(n1769), .A2(n3388), .ZN(n1768) );
  INV_X1 U3145 ( .A(n1364), .ZN(n3889) );
  INV_X1 U3146 ( .A(n3891), .ZN(n3892) );
  NOR2_X1 U3147 ( .A1(n3721), .A2(n3720), .ZN(n3728) );
  INV_X1 U3148 ( .A(n3209), .ZN(n3212) );
  AOI21_X1 U3149 ( .B1(n2757), .B2(n2760), .A(n2758), .ZN(n2718) );
  NOR2_X1 U3150 ( .A1(n2760), .A2(n2757), .ZN(n2717) );
  NAND2_X1 U3153 ( .A1(n2278), .A2(n3193), .ZN(n1736) );
  NAND2_X2 U3154 ( .A1(n2152), .A2(n2050), .ZN(n2151) );
  OAI21_X1 U3155 ( .B1(n2860), .B2(n2847), .A(n2859), .ZN(n2863) );
  NOR3_X4 U3156 ( .A1(n2272), .A2(n2689), .A3(n2316), .ZN(n2315) );
  NAND2_X2 U3157 ( .A1(n1947), .A2(n1953), .ZN(n1513) );
  NAND2_X1 U3159 ( .A1(n1629), .A2(n3237), .ZN(n1520) );
  NAND2_X2 U3160 ( .A1(n1519), .A2(n1518), .ZN(n1521) );
  INV_X2 U3161 ( .A(n1629), .ZN(n1519) );
  OAI21_X1 U3162 ( .B1(n1348), .B2(n2674), .A(n2673), .ZN(n3380) );
  NAND2_X2 U3163 ( .A1(n2204), .A2(n2203), .ZN(n2518) );
  NAND2_X2 U3165 ( .A1(n1524), .A2(n1525), .ZN(\d[27]_BAR ) );
  NAND2_X2 U3166 ( .A1(n1528), .A2(n2007), .ZN(n1530) );
  INV_X1 U3171 ( .A(n3102), .ZN(n3823) );
  NAND2_X2 U3172 ( .A1(a[14]), .A2(n3206), .ZN(n1654) );
  NAND3_X1 U3176 ( .A1(n3920), .A2(n3855), .A3(n3854), .ZN(n3859) );
  INV_X1 U3177 ( .A(n3024), .ZN(n3018) );
  NAND2_X1 U3179 ( .A1(n244), .A2(n2815), .ZN(n1538) );
  NAND2_X1 U3182 ( .A1(n1303), .A2(n3407), .ZN(n2782) );
  NOR2_X1 U3183 ( .A1(n96), .A2(n1303), .ZN(n2169) );
  INV_X1 U3185 ( .A(n2130), .ZN(n2889) );
  NAND2_X1 U3186 ( .A1(n2887), .A2(n2886), .ZN(n2130) );
  INV_X1 U3187 ( .A(n2970), .ZN(n2972) );
  AOI22_X1 U3188 ( .A1(n3132), .A2(n3131), .B1(n3130), .B2(n1487), .ZN(n3182)
         );
  NAND2_X1 U3189 ( .A1(n2852), .A2(n2853), .ZN(n2854) );
  NOR2_X1 U3190 ( .A1(n4008), .A2(n3947), .ZN(n3949) );
  NAND2_X1 U3192 ( .A1(n2026), .A2(n3009), .ZN(n1763) );
  INV_X1 U3193 ( .A(n249), .ZN(n2028) );
  NOR2_X1 U3194 ( .A1(n3177), .A2(n1763), .ZN(n1762) );
  NAND2_X1 U3195 ( .A1(n1350), .A2(n2319), .ZN(n1542) );
  NAND2_X1 U3196 ( .A1(n3450), .A2(n3449), .ZN(n1545) );
  NAND2_X2 U3198 ( .A1(n1545), .A2(n1546), .ZN(n1969) );
  NAND2_X1 U3199 ( .A1(n3436), .A2(n3435), .ZN(n1549) );
  NAND2_X2 U3200 ( .A1(n1549), .A2(n1550), .ZN(n3449) );
  INV_X1 U3201 ( .A(n3436), .ZN(n1547) );
  INV_X1 U3202 ( .A(n3609), .ZN(n3953) );
  NAND2_X1 U3203 ( .A1(n60), .A2(n3609), .ZN(n1894) );
  NAND2_X1 U3205 ( .A1(n1266), .A2(n88), .ZN(n1775) );
  NAND2_X1 U3207 ( .A1(n1507), .A2(n3085), .ZN(n1770) );
  NAND2_X1 U3209 ( .A1(n1261), .A2(a[9]), .ZN(n1977) );
  NAND2_X1 U3210 ( .A1(n1261), .A2(n93), .ZN(n2810) );
  NAND2_X1 U3211 ( .A1(n3427), .A2(a[13]), .ZN(n1814) );
  NAND2_X1 U3212 ( .A1(n1261), .A2(a[20]), .ZN(n1816) );
  NOR2_X1 U3213 ( .A1(n3806), .A2(n3803), .ZN(n3809) );
  NOR2_X1 U3215 ( .A1(n3808), .A2(n3806), .ZN(n1801) );
  NOR2_X2 U3216 ( .A1(n2427), .A2(n2426), .ZN(n2429) );
  NAND2_X4 U3217 ( .A1(n2100), .A2(n4066), .ZN(n3103) );
  AOI22_X1 U3219 ( .A1(n3493), .A2(n1672), .B1(n1968), .B2(n1967), .ZN(n1966)
         );
  NAND2_X2 U3220 ( .A1(n1828), .A2(n1826), .ZN(n3448) );
  INV_X4 U3221 ( .A(n2975), .ZN(n1710) );
  NAND2_X1 U3222 ( .A1(n3794), .A2(n3905), .ZN(n3796) );
  NAND2_X1 U3223 ( .A1(n3804), .A2(n3803), .ZN(n3808) );
  NOR2_X4 U3226 ( .A1(n1774), .A2(n2205), .ZN(\d[29] ) );
  NOR2_X4 U3228 ( .A1(n2180), .A2(n2179), .ZN(n3783) );
  NOR3_X2 U3229 ( .A1(n2074), .A2(n2073), .A3(n2065), .ZN(n3238) );
  NAND3_X2 U3230 ( .A1(n1908), .A2(n1909), .A3(n1906), .ZN(n1568) );
  OAI22_X1 U3231 ( .A1(n3080), .A2(n94), .B1(a[12]), .B2(n1302), .ZN(n2074) );
  NAND2_X1 U3232 ( .A1(n4025), .A2(n2061), .ZN(n4026) );
  AOI21_X1 U3233 ( .B1(n1286), .B2(n2721), .A(n2106), .ZN(n2768) );
  INV_X1 U3235 ( .A(n4026), .ZN(n1572) );
  INV_X4 U3236 ( .A(n2174), .ZN(n1913) );
  NAND2_X2 U3237 ( .A1(n1400), .A2(n1475), .ZN(n1578) );
  INV_X1 U3238 ( .A(n1384), .ZN(n1580) );
  INV_X1 U3239 ( .A(n2029), .ZN(n1583) );
  INV_X2 U3240 ( .A(n1881), .ZN(n1584) );
  AOI21_X1 U3241 ( .B1(n1510), .B2(n4004), .A(n3968), .ZN(n3973) );
  INV_X2 U3242 ( .A(n3799), .ZN(n3814) );
  NAND2_X1 U3243 ( .A1(n3578), .A2(n3577), .ZN(n1586) );
  NOR2_X2 U3246 ( .A1(n3604), .A2(n434), .ZN(n3563) );
  INV_X1 U3247 ( .A(n3679), .ZN(n3676) );
  NAND2_X1 U3249 ( .A1(n2147), .A2(n675), .ZN(n1593) );
  NAND2_X1 U3250 ( .A1(n3721), .A2(n3720), .ZN(n3716) );
  INV_X2 U3251 ( .A(n3785), .ZN(n3797) );
  INV_X1 U3253 ( .A(n2066), .ZN(n3968) );
  INV_X4 U3255 ( .A(b[8]), .ZN(n1596) );
  NOR2_X1 U3256 ( .A1(n1392), .A2(n3793), .ZN(n3750) );
  OAI21_X2 U3258 ( .B1(n1471), .B2(n3603), .A(n1540), .ZN(n1601) );
  NAND2_X1 U3260 ( .A1(n3328), .A2(n2084), .ZN(n3209) );
  NAND2_X1 U3261 ( .A1(n45), .A2(n1449), .ZN(n2459) );
  OAI21_X1 U3263 ( .B1(n1244), .B2(n3294), .A(n3293), .ZN(n1640) );
  NAND2_X1 U3264 ( .A1(n1517), .A2(n1208), .ZN(n3279) );
  NAND2_X1 U3267 ( .A1(n2980), .A2(n2355), .ZN(n1858) );
  INV_X1 U3268 ( .A(n1498), .ZN(n3756) );
  INV_X4 U3269 ( .A(n3034), .ZN(n1705) );
  NAND2_X1 U3270 ( .A1(n3203), .A2(a[3]), .ZN(n3014) );
  NOR2_X1 U3271 ( .A1(n3203), .A2(n3128), .ZN(n2171) );
  NAND2_X1 U3272 ( .A1(n3203), .A2(n56), .ZN(n2379) );
  NOR2_X1 U3273 ( .A1(n3203), .A2(n3202), .ZN(n2073) );
  MUX2_X2 U3275 ( .A(n1361), .B(n3203), .S(n3468), .Z(n2867) );
  AOI22_X1 U3276 ( .A1(n3996), .A2(n1892), .B1(n4019), .B2(n3990), .ZN(n3992)
         );
  NOR2_X1 U3277 ( .A1(n1453), .A2(n3505), .ZN(n3508) );
  NOR2_X1 U3278 ( .A1(n3514), .A2(n1453), .ZN(n3520) );
  INV_X1 U3279 ( .A(n3293), .ZN(n2126) );
  NOR3_X1 U3280 ( .A1(n3828), .A2(n3827), .A3(n3907), .ZN(n3835) );
  NAND2_X1 U3281 ( .A1(n3371), .A2(n2088), .ZN(n2152) );
  NAND2_X1 U3282 ( .A1(n1927), .A2(n4010), .ZN(n3964) );
  INV_X1 U3284 ( .A(n2481), .ZN(n2479) );
  INV_X4 U3286 ( .A(n1928), .ZN(n1863) );
  NAND2_X1 U3288 ( .A1(n3034), .A2(n2079), .ZN(n2078) );
  NAND2_X1 U3289 ( .A1(n3034), .A2(n2077), .ZN(n1982) );
  NOR2_X1 U3290 ( .A1(n1303), .A2(a[8]), .ZN(n2832) );
  NOR2_X1 U3292 ( .A1(n3328), .A2(a[8]), .ZN(n1993) );
  XNOR2_X1 U3293 ( .A(a[8]), .B(n2200), .ZN(n3017) );
  NAND3_X1 U3294 ( .A1(n3067), .A2(a[8]), .A3(n2506), .ZN(n3068) );
  OAI21_X1 U3295 ( .B1(n3517), .B2(n2356), .A(n916), .ZN(n3518) );
  NAND2_X1 U3296 ( .A1(n2356), .A2(n1261), .ZN(n2324) );
  NAND2_X1 U3297 ( .A1(n2356), .A2(n3453), .ZN(n1974) );
  XNOR2_X1 U3298 ( .A(n92), .B(a[25]), .ZN(n3643) );
  NAND3_X1 U3299 ( .A1(n3010), .A2(n2907), .A3(n2356), .ZN(n1919) );
  AOI21_X1 U3300 ( .B1(n249), .B2(n3538), .A(n3010), .ZN(n2999) );
  INV_X4 U3302 ( .A(n1836), .ZN(n1837) );
  NAND2_X2 U3304 ( .A1(n1639), .A2(n1623), .ZN(n4009) );
  NAND2_X2 U3305 ( .A1(n1617), .A2(n1622), .ZN(n1621) );
  INV_X4 U3307 ( .A(n1729), .ZN(n3052) );
  OAI22_X2 U3308 ( .A1(n2144), .A2(n92), .B1(n2143), .B2(n2997), .ZN(n2954) );
  INV_X4 U3309 ( .A(n3013), .ZN(n3054) );
  INV_X2 U3310 ( .A(n3278), .ZN(n1955) );
  OAI22_X2 U3311 ( .A1(n3763), .A2(n1677), .B1(n3761), .B2(n3762), .ZN(n1973)
         );
  NAND2_X2 U3312 ( .A1(n1676), .A2(n1675), .ZN(n3763) );
  AOI22_X2 U3314 ( .A1(n2982), .A2(n1687), .B1(n1859), .B2(n3589), .ZN(n2559)
         );
  INV_X4 U3315 ( .A(n2936), .ZN(n2226) );
  OAI21_X2 U3316 ( .B1(n1331), .B2(n2138), .A(n1635), .ZN(n2135) );
  NAND3_X2 U3317 ( .A1(n1779), .A2(n1707), .A3(n2380), .ZN(n2342) );
  NAND2_X2 U3318 ( .A1(n1641), .A2(n471), .ZN(n1644) );
  NAND2_X2 U3319 ( .A1(n1643), .A2(n1642), .ZN(n1641) );
  NAND2_X2 U3320 ( .A1(n1777), .A2(n3355), .ZN(n1642) );
  NAND2_X2 U3321 ( .A1(n1645), .A2(n444), .ZN(n1931) );
  OAI21_X1 U3322 ( .B1(n3495), .B2(n1645), .A(n2476), .ZN(n2463) );
  INV_X4 U3323 ( .A(n3026), .ZN(n1645) );
  INV_X2 U3324 ( .A(n1928), .ZN(n1862) );
  OAI21_X2 U3326 ( .B1(n3924), .B2(n3693), .A(n1648), .ZN(n3694) );
  NOR3_X2 U3327 ( .A1(n3692), .A2(n3690), .A3(n3691), .ZN(n1648) );
  INV_X4 U3329 ( .A(n2830), .ZN(n3839) );
  BUF_X4 U3330 ( .A(n3431), .Z(n1649) );
  NOR2_X2 U3332 ( .A1(n3777), .A2(n1925), .ZN(n1650) );
  BUF_X4 U3333 ( .A(b[7]), .Z(n1651) );
  NAND2_X2 U3335 ( .A1(n1449), .A2(n2438), .ZN(n1653) );
  NAND3_X2 U3336 ( .A1(n2035), .A2(n2036), .A3(n2037), .ZN(n3168) );
  NOR3_X2 U3337 ( .A1(n4046), .A2(n2273), .A3(n451), .ZN(n1753) );
  NAND2_X2 U3339 ( .A1(n2096), .A2(n2810), .ZN(n2095) );
  NAND3_X2 U3341 ( .A1(n1656), .A2(n3697), .A3(n3696), .ZN(\d[36] ) );
  INV_X2 U3342 ( .A(n2954), .ZN(n2142) );
  INV_X1 U3343 ( .A(n1857), .ZN(n1773) );
  NAND2_X2 U3344 ( .A1(n2654), .A2(a[1]), .ZN(n1658) );
  AOI21_X2 U3345 ( .B1(n3061), .B2(n3062), .A(n3059), .ZN(n3049) );
  NOR2_X2 U3346 ( .A1(n1664), .A2(n1662), .ZN(n1677) );
  NAND2_X2 U3347 ( .A1(n1663), .A2(n3762), .ZN(n1662) );
  INV_X2 U3348 ( .A(n3555), .ZN(n1663) );
  NAND3_X2 U3349 ( .A1(n1669), .A2(n1668), .A3(n1667), .ZN(n1676) );
  XNOR2_X2 U3350 ( .A(n3540), .B(n3539), .ZN(n1668) );
  NOR2_X2 U3352 ( .A1(n1671), .A2(n3541), .ZN(n1670) );
  INV_X2 U3353 ( .A(n3524), .ZN(n1671) );
  BUF_X4 U3354 ( .A(n3542), .Z(n1672) );
  NAND2_X2 U3355 ( .A1(n1674), .A2(n1673), .ZN(n1675) );
  NAND2_X2 U3356 ( .A1(n1679), .A2(n1678), .ZN(n3761) );
  NAND2_X2 U3357 ( .A1(n1396), .A2(n464), .ZN(n1678) );
  NAND2_X2 U3359 ( .A1(n2361), .A2(n2856), .ZN(n1682) );
  AOI21_X1 U3360 ( .B1(n1684), .B2(n2945), .A(n2944), .ZN(n3172) );
  NAND2_X2 U3361 ( .A1(n2436), .A2(n2437), .ZN(n1689) );
  NAND2_X2 U3364 ( .A1(n2396), .A2(n1316), .ZN(n1772) );
  NAND2_X2 U3365 ( .A1(n1696), .A2(n3242), .ZN(n1695) );
  XNOR2_X2 U3366 ( .A(n1706), .B(n2924), .ZN(n2271) );
  OAI22_X2 U3367 ( .A1(n1589), .A2(n1708), .B1(n3101), .B2(n68), .ZN(n1937) );
  NAND2_X2 U3368 ( .A1(n1710), .A2(n2976), .ZN(n3086) );
  INV_X4 U3369 ( .A(n3065), .ZN(n1890) );
  NOR2_X2 U3371 ( .A1(n3888), .A2(n1243), .ZN(n3886) );
  NAND2_X1 U3373 ( .A1(n3472), .A2(n98), .ZN(n1715) );
  NAND2_X1 U3376 ( .A1(n2438), .A2(n3455), .ZN(n2387) );
  NAND2_X1 U3377 ( .A1(n1016), .A2(n3016), .ZN(n2796) );
  MUX2_X2 U3378 ( .A(n1016), .B(n3472), .S(a[8]), .Z(n2996) );
  MUX2_X2 U3379 ( .A(n1016), .B(n3472), .S(a[11]), .Z(n2865) );
  MUX2_X2 U3380 ( .A(n1016), .B(n3472), .S(a[10]), .Z(n2895) );
  NAND2_X2 U3381 ( .A1(n1723), .A2(n1722), .ZN(n2855) );
  NAND2_X2 U3382 ( .A1(n1721), .A2(n3534), .ZN(n1996) );
  OAI21_X2 U3386 ( .B1(n3054), .B2(n3058), .A(n3012), .ZN(n3061) );
  OAI22_X2 U3389 ( .A1(n3001), .A2(n1705), .B1(n2999), .B2(n3000), .ZN(n3051)
         );
  NAND2_X4 U3390 ( .A1(n2740), .A2(n1735), .ZN(n3080) );
  NAND2_X2 U3391 ( .A1(n3515), .A2(n1735), .ZN(n3332) );
  NAND2_X2 U3392 ( .A1(n1736), .A2(n3164), .ZN(n2234) );
  NAND2_X2 U3393 ( .A1(n1737), .A2(n2129), .ZN(n1983) );
  INV_X2 U3394 ( .A(n1743), .ZN(n1742) );
  NOR2_X2 U3395 ( .A1(n1744), .A2(n2232), .ZN(n1743) );
  NOR2_X1 U3396 ( .A1(n1745), .A2(n3909), .ZN(n3912) );
  AOI21_X2 U3398 ( .B1(n2526), .B2(n2208), .A(n2565), .ZN(n2527) );
  OAI21_X2 U3399 ( .B1(n1748), .B2(n1747), .A(n1746), .ZN(n3450) );
  XNOR2_X2 U3400 ( .A(n1749), .B(n3452), .ZN(n3487) );
  INV_X2 U3401 ( .A(n1751), .ZN(n2988) );
  NAND2_X2 U3402 ( .A1(n2830), .A2(n1752), .ZN(n1751) );
  NAND2_X2 U3403 ( .A1(n1756), .A2(n1753), .ZN(n2852) );
  NOR2_X4 U3405 ( .A1(n1207), .A2(n3095), .ZN(n3825) );
  NAND2_X2 U3406 ( .A1(n2889), .A2(n1751), .ZN(n1760) );
  INV_X4 U3407 ( .A(n3020), .ZN(n1830) );
  NOR2_X2 U3408 ( .A1(n2390), .A2(n1084), .ZN(n2827) );
  NAND2_X2 U3409 ( .A1(n3327), .A2(n3326), .ZN(n1769) );
  NAND2_X2 U3410 ( .A1(n1379), .A2(n1770), .ZN(n2100) );
  NAND3_X2 U3411 ( .A1(n3557), .A2(n1408), .A3(n2012), .ZN(n1771) );
  INV_X2 U3412 ( .A(n4021), .ZN(n1804) );
  NAND3_X2 U3413 ( .A1(n3943), .A2(n3942), .A3(n3941), .ZN(n1774) );
  INV_X4 U3414 ( .A(n3206), .ZN(n2070) );
  NAND2_X2 U3415 ( .A1(n3522), .A2(n2941), .ZN(n1776) );
  BUF_X4 U3416 ( .A(n3353), .Z(n1777) );
  AOI21_X2 U3420 ( .B1(n1982), .B2(n4057), .A(n2997), .ZN(n1780) );
  AOI21_X2 U3422 ( .B1(n1981), .B2(n2123), .A(n92), .ZN(n1783) );
  BUF_X4 U3423 ( .A(a[4]), .Z(n1784) );
  INV_X2 U3424 ( .A(n3199), .ZN(n1852) );
  BUF_X4 U3425 ( .A(n3910), .Z(n1787) );
  BUF_X4 U3426 ( .A(n3164), .Z(n1788) );
  OAI21_X2 U3430 ( .B1(n3807), .B2(n1802), .A(n1799), .ZN(\d[12]_BAR ) );
  NOR2_X2 U3431 ( .A1(n1801), .A2(n4060), .ZN(n1799) );
  NAND2_X2 U3433 ( .A1(n1272), .A2(n1445), .ZN(n1803) );
  BUF_X4 U3434 ( .A(n3810), .Z(n2320) );
  NAND3_X1 U3435 ( .A1(n3999), .A2(n4070), .A3(n4015), .ZN(n4000) );
  INV_X8 U3436 ( .A(n2359), .ZN(n3431) );
  NAND2_X4 U3437 ( .A1(n1898), .A2(n3065), .ZN(n2359) );
  NAND3_X2 U3438 ( .A1(n1808), .A2(n3992), .A3(n3991), .ZN(n4002) );
  AOI21_X2 U3439 ( .B1(n2226), .B2(n2937), .A(n2377), .ZN(n3981) );
  NAND2_X4 U3440 ( .A1(n3129), .A2(n1818), .ZN(n3310) );
  NAND3_X1 U3442 ( .A1(n1487), .A2(n1818), .A3(n3202), .ZN(n1815) );
  NAND2_X2 U3443 ( .A1(n1817), .A2(n1816), .ZN(n2402) );
  NAND3_X1 U3444 ( .A1(n1487), .A2(n1818), .A3(n3109), .ZN(n1817) );
  INV_X4 U3445 ( .A(n3127), .ZN(n1818) );
  NAND2_X2 U3446 ( .A1(n85), .A2(n2228), .ZN(n2096) );
  MUX2_X2 U3447 ( .A(n85), .B(n1261), .S(a[21]), .Z(n2427) );
  MUX2_X2 U3448 ( .A(n85), .B(n1261), .S(a[12]), .Z(n2843) );
  MUX2_X2 U3449 ( .A(n85), .B(n1261), .S(a[19]), .Z(n2408) );
  NOR2_X2 U3451 ( .A1(n2516), .A2(n2441), .ZN(n1822) );
  NAND2_X2 U3452 ( .A1(n1825), .A2(n16), .ZN(n2522) );
  NAND3_X2 U3453 ( .A1(n1827), .A2(n3783), .A3(n4067), .ZN(n1826) );
  INV_X2 U3454 ( .A(n1576), .ZN(n1827) );
  NAND2_X2 U3455 ( .A1(n2173), .A2(n2172), .ZN(n3441) );
  INV_X8 U3457 ( .A(b[13]), .ZN(n2924) );
  INV_X2 U3459 ( .A(n2924), .ZN(n1836) );
  OR2_X4 U3460 ( .A1(n2924), .A2(b[14]), .ZN(n1835) );
  NAND2_X2 U3461 ( .A1(n3260), .A2(n3259), .ZN(n1838) );
  NAND2_X2 U3463 ( .A1(n1377), .A2(n3413), .ZN(n2781) );
  INV_X1 U3464 ( .A(n2946), .ZN(n1839) );
  INV_X2 U3465 ( .A(n2933), .ZN(n1841) );
  INV_X2 U3466 ( .A(n3360), .ZN(n1843) );
  NOR2_X2 U3467 ( .A1(n1464), .A2(n1844), .ZN(n3360) );
  INV_X8 U3468 ( .A(n1845), .ZN(n3328) );
  NAND2_X2 U3469 ( .A1(n2348), .A2(n2346), .ZN(n2910) );
  NAND2_X4 U3470 ( .A1(n1846), .A2(n3618), .ZN(n3920) );
  NAND2_X2 U3471 ( .A1(n3611), .A2(n1848), .ZN(n1847) );
  NOR2_X4 U3472 ( .A1(n1849), .A2(n3675), .ZN(n3618) );
  NAND2_X4 U3473 ( .A1(n3707), .A2(n3711), .ZN(n3675) );
  NAND2_X2 U3474 ( .A1(n3578), .A2(n3577), .ZN(n3707) );
  NOR2_X2 U3475 ( .A1(n3720), .A2(n1850), .ZN(n1849) );
  NOR2_X4 U3476 ( .A1(n3577), .A2(n3578), .ZN(n3720) );
  NAND2_X2 U3477 ( .A1(n1853), .A2(n3199), .ZN(n3133) );
  NAND2_X2 U3478 ( .A1(n2110), .A2(n2107), .ZN(n2721) );
  NAND2_X2 U3479 ( .A1(n1864), .A2(n1856), .ZN(n2188) );
  NAND2_X2 U3480 ( .A1(n2981), .A2(n1858), .ZN(n2113) );
  NAND2_X2 U3481 ( .A1(n1861), .A2(n1860), .ZN(n2985) );
  NOR2_X2 U3482 ( .A1(n2876), .A2(n2877), .ZN(n1874) );
  INV_X2 U3483 ( .A(n3103), .ZN(n3757) );
  INV_X2 U3485 ( .A(n2721), .ZN(n1875) );
  INV_X8 U3486 ( .A(n2165), .ZN(n3177) );
  INV_X4 U3488 ( .A(n3186), .ZN(n3180) );
  NAND2_X2 U3490 ( .A1(n2362), .A2(n2855), .ZN(n2361) );
  NAND3_X2 U3491 ( .A1(n4047), .A2(n1996), .A3(n1994), .ZN(n2362) );
  XNOR2_X1 U3494 ( .A(n2924), .B(a[10]), .ZN(n3143) );
  AOI22_X2 U3495 ( .A1(n3140), .A2(n3010), .B1(n3141), .B2(n1837), .ZN(n3142)
         );
  NAND2_X1 U3498 ( .A1(n1889), .A2(n1898), .ZN(n1888) );
  BUF_X4 U3499 ( .A(n3933), .Z(n1892) );
  NAND2_X2 U3500 ( .A1(n2310), .A2(n2566), .ZN(n2309) );
  NOR2_X4 U3501 ( .A1(n3872), .A2(n3871), .ZN(n3929) );
  NOR3_X2 U3502 ( .A1(n1897), .A2(n4010), .A3(n1938), .ZN(n3871) );
  AOI21_X2 U3503 ( .B1(n1409), .B2(n3609), .A(n3720), .ZN(n1895) );
  INV_X1 U3504 ( .A(n3606), .ZN(n1896) );
  NAND2_X2 U3505 ( .A1(n3496), .A2(n4155), .ZN(n3500) );
  INV_X2 U3506 ( .A(n2331), .ZN(n1901) );
  INV_X2 U3507 ( .A(n1911), .ZN(n2357) );
  NAND2_X2 U3508 ( .A1(n1907), .A2(n4156), .ZN(n1906) );
  INV_X4 U3509 ( .A(b[1]), .ZN(n2556) );
  INV_X2 U3514 ( .A(n964), .ZN(n1925) );
  NOR2_X1 U3515 ( .A1(n3954), .A2(n1497), .ZN(n1927) );
  NAND2_X2 U3517 ( .A1(n1930), .A2(n4049), .ZN(n2177) );
  INV_X4 U3518 ( .A(n2072), .ZN(n2856) );
  INV_X4 U3519 ( .A(n1898), .ZN(n3026) );
  NAND2_X2 U3521 ( .A1(n1935), .A2(n1934), .ZN(n1936) );
  INV_X2 U3522 ( .A(n1483), .ZN(n3285) );
  INV_X4 U3523 ( .A(n2980), .ZN(n2737) );
  NOR2_X4 U3524 ( .A1(n1943), .A2(n2623), .ZN(n2674) );
  INV_X1 U3525 ( .A(n1578), .ZN(n3815) );
  NAND3_X1 U3526 ( .A1(n3799), .A2(n3785), .A3(n1578), .ZN(n2089) );
  NAND2_X1 U3527 ( .A1(n3813), .A2(n1578), .ZN(n3801) );
  NAND3_X2 U3529 ( .A1(n1952), .A2(n1949), .A3(n1948), .ZN(n3278) );
  NAND2_X2 U3532 ( .A1(n95), .A2(n85), .ZN(n2325) );
  MUX2_X2 U3533 ( .A(n85), .B(n1261), .S(n3538), .Z(n3428) );
  MUX2_X2 U3534 ( .A(n85), .B(n1261), .S(a[1]), .Z(n3393) );
  MUX2_X2 U3535 ( .A(n85), .B(n1261), .S(n205), .Z(n3002) );
  NAND2_X2 U3536 ( .A1(n2241), .A2(n2240), .ZN(n2916) );
  NAND2_X2 U3538 ( .A1(n3480), .A2(n3487), .ZN(n1968) );
  NOR2_X2 U3539 ( .A1(n3769), .A2(n3491), .ZN(n3766) );
  NAND2_X2 U3540 ( .A1(n1975), .A2(n1974), .ZN(n3457) );
  MUX2_X2 U3541 ( .A(n3200), .B(n3453), .S(a[3]), .Z(n3406) );
  MUX2_X2 U3542 ( .A(n1976), .B(n3453), .S(a[8]), .Z(n3082) );
  INV_X4 U3543 ( .A(n3289), .ZN(n2128) );
  NOR2_X2 U3544 ( .A1(n1804), .A2(n3661), .ZN(n3662) );
  NAND2_X2 U3545 ( .A1(n3609), .A2(n3956), .ZN(n2248) );
  NAND2_X2 U3546 ( .A1(n1990), .A2(n2191), .ZN(n3609) );
  XNOR2_X2 U3547 ( .A(n2462), .B(n1998), .ZN(n1997) );
  AOI21_X2 U3548 ( .B1(n3143), .B2(n313), .A(n3142), .ZN(n3186) );
  INV_X4 U3549 ( .A(n3989), .ZN(n1999) );
  NOR2_X2 U3550 ( .A1(n2002), .A2(n2001), .ZN(n3989) );
  NOR2_X2 U3551 ( .A1(n2008), .A2(n2327), .ZN(n2006) );
  NOR2_X4 U3552 ( .A1(n2010), .A2(n2357), .ZN(n3298) );
  INV_X4 U3554 ( .A(n3208), .ZN(n3113) );
  NAND2_X2 U3555 ( .A1(n2453), .A2(n476), .ZN(n2455) );
  NAND2_X2 U3556 ( .A1(n2288), .A2(n2014), .ZN(n2289) );
  NAND2_X2 U3557 ( .A1(n2017), .A2(n2016), .ZN(n2015) );
  INV_X2 U3558 ( .A(n2923), .ZN(n2016) );
  INV_X2 U3559 ( .A(n2223), .ZN(n2017) );
  NAND3_X2 U3560 ( .A1(n1542), .A2(n3557), .A3(n3556), .ZN(n3810) );
  NOR2_X2 U3561 ( .A1(n2019), .A2(n3535), .ZN(n3536) );
  INV_X1 U3562 ( .A(n3496), .ZN(n2019) );
  NAND3_X1 U3563 ( .A1(n313), .A2(n2997), .A3(n96), .ZN(n2023) );
  MUX2_X2 U3566 ( .A(n2980), .B(n2022), .S(a[23]), .Z(n2683) );
  NAND2_X2 U3568 ( .A1(n2113), .A2(n1773), .ZN(n2995) );
  NAND3_X2 U3570 ( .A1(n2034), .A2(n2033), .A3(n2032), .ZN(n2035) );
  NOR2_X2 U3571 ( .A1(n1285), .A2(n2081), .ZN(n2034) );
  INV_X4 U3572 ( .A(n2688), .ZN(n2272) );
  NAND2_X2 U3573 ( .A1(b[8]), .A2(b[7]), .ZN(n2688) );
  NAND3_X1 U3574 ( .A1(n2045), .A2(n3177), .A3(n1836), .ZN(n2044) );
  AOI21_X2 U3575 ( .B1(n1914), .B2(n2893), .A(n1280), .ZN(n2881) );
  NAND2_X2 U3576 ( .A1(n2215), .A2(n1166), .ZN(n2048) );
  NAND2_X2 U3578 ( .A1(n2178), .A2(n2937), .ZN(n2055) );
  NOR2_X2 U3579 ( .A1(n2058), .A2(a[9]), .ZN(n2822) );
  MUX2_X2 U3584 ( .A(n86), .B(n2058), .S(n2407), .Z(n2424) );
  MUX2_X2 U3585 ( .A(n155), .B(n2058), .S(n3217), .Z(n2591) );
  INV_X4 U3586 ( .A(n3328), .ZN(n2058) );
  OAI22_X2 U3587 ( .A1(n3625), .A2(n3626), .B1(n3624), .B2(n3623), .ZN(
        \d[37]_BAR ) );
  OAI22_X2 U3589 ( .A1(n2062), .A2(n2060), .B1(n3701), .B2(n2061), .ZN(n3703)
         );
  NAND2_X2 U3590 ( .A1(n3701), .A2(n2061), .ZN(n2060) );
  BUF_X4 U3591 ( .A(n4003), .Z(n2066) );
  NOR2_X2 U3592 ( .A1(n2485), .A2(n2484), .ZN(n2503) );
  NAND2_X4 U3593 ( .A1(b[9]), .A2(b[10]), .ZN(n2741) );
  INV_X8 U3594 ( .A(b[5]), .ZN(n2785) );
  NOR2_X2 U3596 ( .A1(n3571), .A2(n3570), .ZN(n3910) );
  INV_X4 U3597 ( .A(n1362), .ZN(n3145) );
  AOI21_X2 U3598 ( .B1(n1238), .B2(n3157), .A(n3156), .ZN(n2081) );
  INV_X8 U3599 ( .A(n3003), .ZN(n3329) );
  INV_X8 U3600 ( .A(n2315), .ZN(n3323) );
  AOI21_X2 U3605 ( .B1(n836), .B2(n4016), .A(n4014), .ZN(\d[26] ) );
  NOR2_X2 U3607 ( .A1(n2353), .A2(n2094), .ZN(n2093) );
  INV_X1 U3608 ( .A(n2859), .ZN(n2813) );
  NOR2_X2 U3610 ( .A1(n2110), .A2(n2107), .ZN(n2106) );
  NAND2_X1 U3611 ( .A1(n1361), .A2(n3139), .ZN(n2378) );
  NAND2_X1 U3612 ( .A1(n84), .A2(n3534), .ZN(n3015) );
  MUX2_X2 U3613 ( .A(n3203), .B(n3080), .S(n2438), .Z(n2554) );
  MUX2_X2 U3614 ( .A(n3203), .B(n1361), .S(n2613), .Z(n2681) );
  NOR2_X2 U3615 ( .A1(n3104), .A2(n3103), .ZN(n3883) );
  INV_X4 U3616 ( .A(n857), .ZN(n2199) );
  NAND2_X1 U3618 ( .A1(n4074), .A2(n1224), .ZN(n2873) );
  NOR2_X1 U3619 ( .A1(n4074), .A2(n1224), .ZN(n2874) );
  NAND2_X1 U3620 ( .A1(n3186), .A2(n2120), .ZN(n3156) );
  NOR2_X2 U3623 ( .A1(n2248), .A2(n3994), .ZN(n2129) );
  NAND3_X2 U3626 ( .A1(n1349), .A2(n1219), .A3(n2136), .ZN(n2134) );
  INV_X2 U3627 ( .A(n1766), .ZN(n3513) );
  NOR2_X2 U3628 ( .A1(n2223), .A2(n2923), .ZN(n2953) );
  AOI22_X2 U3629 ( .A1(n3373), .A2(n446), .B1(n1324), .B2(n1310), .ZN(n2148)
         );
  NOR2_X1 U3632 ( .A1(n3016), .A2(n2316), .ZN(n2347) );
  XNOR2_X1 U3633 ( .A(n2316), .B(n2412), .ZN(n2413) );
  NOR2_X2 U3634 ( .A1(n2377), .A2(n2226), .ZN(n2178) );
  AOI22_X2 U3636 ( .A1(n3435), .A2(n3395), .B1(n2182), .B2(n3394), .ZN(n3419)
         );
  INV_X4 U3637 ( .A(n2185), .ZN(n3170) );
  NAND2_X2 U3639 ( .A1(n2190), .A2(n18), .ZN(n2189) );
  INV_X4 U3640 ( .A(b[2]), .ZN(n3066) );
  NOR2_X2 U3641 ( .A1(n1400), .A2(n1475), .ZN(n3817) );
  INV_X4 U3642 ( .A(n3027), .ZN(n2200) );
  NAND2_X2 U3643 ( .A1(n3453), .A2(a[22]), .ZN(n2203) );
  NAND2_X2 U3644 ( .A1(n3946), .A2(n3944), .ZN(n2206) );
  INV_X2 U3645 ( .A(n3117), .ZN(n3116) );
  NAND2_X2 U3646 ( .A1(n2213), .A2(n2210), .ZN(n3117) );
  NOR2_X2 U3647 ( .A1(n2212), .A2(n2211), .ZN(n2210) );
  NOR2_X1 U3648 ( .A1(n3328), .A2(n94), .ZN(n2211) );
  NOR2_X1 U3649 ( .A1(n2084), .A2(n3202), .ZN(n2212) );
  NOR2_X4 U3651 ( .A1(n3129), .A2(n3125), .ZN(n3427) );
  NAND2_X2 U3652 ( .A1(n2225), .A2(n2224), .ZN(n2223) );
  BUF_X4 U3653 ( .A(n3162), .Z(n2230) );
  XNOR2_X1 U3654 ( .A(n1323), .B(n2026), .ZN(n3073) );
  XNOR2_X1 U3655 ( .A(n1323), .B(n2239), .ZN(n3211) );
  XNOR2_X1 U3656 ( .A(n1323), .B(a[7]), .ZN(n2885) );
  NAND3_X2 U3657 ( .A1(n2831), .A2(n4034), .A3(n2243), .ZN(n2242) );
  AOI21_X2 U3658 ( .B1(n2601), .B2(n1496), .A(n2250), .ZN(n2249) );
  INV_X2 U3659 ( .A(n2600), .ZN(n2250) );
  NAND2_X2 U3662 ( .A1(n2256), .A2(n2255), .ZN(n2254) );
  INV_X2 U3663 ( .A(n2463), .ZN(n2255) );
  NAND2_X2 U3664 ( .A1(n733), .A2(n2478), .ZN(n2256) );
  NOR2_X2 U3665 ( .A1(n2505), .A2(n2259), .ZN(n2507) );
  NAND2_X2 U3666 ( .A1(n1330), .A2(n2260), .ZN(n2259) );
  AOI21_X2 U3667 ( .B1(n378), .B2(n1631), .A(n3269), .ZN(n3268) );
  XNOR2_X2 U3670 ( .A(n2264), .B(n3908), .ZN(\d[17] ) );
  NOR2_X2 U3671 ( .A1(n3905), .A2(n3904), .ZN(n2264) );
  NAND2_X1 U3672 ( .A1(n1303), .A2(n100), .ZN(n2270) );
  NAND2_X1 U3673 ( .A1(n3823), .A2(n1418), .ZN(n3830) );
  NOR2_X1 U3674 ( .A1(n3328), .A2(a[7]), .ZN(n2273) );
  NAND2_X2 U3675 ( .A1(n2951), .A2(n3145), .ZN(n2278) );
  NOR2_X2 U3677 ( .A1(n2956), .A2(n2959), .ZN(n3160) );
  XNOR2_X1 U3679 ( .A(n1257), .B(n3981), .ZN(n3983) );
  INV_X2 U3680 ( .A(n2289), .ZN(n3963) );
  NOR2_X1 U3681 ( .A1(a[3]), .A2(n2359), .ZN(n2291) );
  INV_X2 U3682 ( .A(n2872), .ZN(n2300) );
  INV_X2 U3683 ( .A(n3729), .ZN(n2308) );
  INV_X8 U3686 ( .A(n2399), .ZN(n3204) );
  NAND2_X4 U3687 ( .A1(n2742), .A2(n2741), .ZN(n3203) );
  INV_X8 U3688 ( .A(n2423), .ZN(n2316) );
  NAND2_X1 U3689 ( .A1(n2315), .A2(a[17]), .ZN(n2389) );
  AOI21_X2 U3691 ( .B1(n2320), .B2(n3786), .A(n3797), .ZN(n3790) );
  NOR2_X2 U3692 ( .A1(n3403), .A2(n3402), .ZN(n2323) );
  NAND2_X2 U3693 ( .A1(n2325), .A2(n2324), .ZN(n3402) );
  NAND3_X2 U3694 ( .A1(n1365), .A2(n3282), .A3(n2328), .ZN(n2326) );
  AOI21_X2 U3695 ( .B1(n1365), .B2(n3282), .A(n2328), .ZN(n2327) );
  NAND3_X2 U3696 ( .A1(n2506), .A2(n2334), .A3(n2333), .ZN(n2332) );
  NAND2_X2 U3698 ( .A1(n3105), .A2(n1322), .ZN(n3891) );
  NAND2_X2 U3699 ( .A1(n1318), .A2(n3883), .ZN(n2341) );
  NOR2_X2 U3700 ( .A1(n3906), .A2(n3825), .ZN(n2343) );
  INV_X2 U3701 ( .A(n3046), .ZN(n2345) );
  INV_X8 U3702 ( .A(b[7]), .ZN(n3027) );
  AOI22_X1 U3703 ( .A1(n3003), .A2(n3016), .B1(n3392), .B2(n2347), .ZN(n2346)
         );
  INV_X4 U3705 ( .A(n3328), .ZN(n2354) );
  INV_X8 U3706 ( .A(n2355), .ZN(n2356) );
  NAND2_X2 U3708 ( .A1(n2367), .A2(n2365), .ZN(n2364) );
  NAND2_X2 U3710 ( .A1(n2369), .A2(n3950), .ZN(n3951) );
  INV_X2 U3711 ( .A(n3948), .ZN(n2369) );
  NAND2_X2 U3712 ( .A1(n2375), .A2(n2370), .ZN(n2374) );
  NAND2_X2 U3713 ( .A1(n2375), .A2(n2373), .ZN(n2846) );
  NAND2_X2 U3715 ( .A1(n2379), .A2(n2378), .ZN(n2835) );
  NAND2_X2 U3717 ( .A1(n3561), .A2(n3100), .ZN(n2380) );
  NAND2_X1 U3718 ( .A1(n1202), .A2(n4011), .ZN(n2381) );
  OAI21_X1 U3720 ( .B1(n2786), .B2(n1245), .A(n2506), .ZN(n2787) );
  XOR2_X1 U3721 ( .A(n25), .B(n3760), .Z(n3771) );
  NAND2_X1 U3722 ( .A1(n4019), .A2(n951), .ZN(n4020) );
  NAND2_X1 U3723 ( .A1(n3024), .A2(n3039), .ZN(n3019) );
  NAND2_X1 U3725 ( .A1(a[13]), .A2(n2145), .ZN(n2798) );
  NOR2_X1 U3726 ( .A1(n3016), .A2(n3498), .ZN(n2882) );
  XNOR2_X1 U3727 ( .A(a[21]), .B(n3122), .ZN(n2516) );
  INV_X1 U3728 ( .A(n3057), .ZN(n3012) );
  NAND3_X1 U3729 ( .A1(n3510), .A2(n2355), .A3(n1752), .ZN(n3511) );
  NAND3_X1 U3730 ( .A1(n3062), .A2(n3060), .A3(n1290), .ZN(n3063) );
  INV_X1 U3731 ( .A(n3259), .ZN(n3261) );
  INV_X1 U3732 ( .A(n3583), .ZN(n3584) );
  OAI21_X1 U3733 ( .B1(n2745), .B2(n2748), .A(n2746), .ZN(n3874) );
  INV_X1 U3734 ( .A(n1586), .ZN(n3708) );
  XNOR2_X1 U3735 ( .A(n3646), .B(n3645), .ZN(n3598) );
  NAND2_X1 U3737 ( .A1(n3483), .A2(n3492), .ZN(n3489) );
  NAND2_X1 U3738 ( .A1(n3450), .A2(n3449), .ZN(n3438) );
  NOR3_X1 U3739 ( .A1(n3766), .A2(n3765), .A3(n3764), .ZN(n3767) );
  NOR3_X1 U3740 ( .A1(n4031), .A2(n3619), .A3(n3621), .ZN(n3601) );
  XNOR2_X1 U3741 ( .A(n185), .B(n1271), .ZN(n3778) );
  XNOR2_X1 U3742 ( .A(n3781), .B(n3782), .ZN(\d[9]_BAR ) );
  BUF_X4 U3743 ( .A(b[11]), .Z(n2740) );
  BUF_X4 U3744 ( .A(b[10]), .Z(n2412) );
  INV_X4 U3745 ( .A(n1448), .ZN(n2399) );
  INV_X4 U3746 ( .A(a[16]), .ZN(n2400) );
  INV_X4 U3748 ( .A(b[6]), .ZN(n3129) );
  NAND2_X2 U3749 ( .A1(n2785), .A2(b[7]), .ZN(n3127) );
  INV_X4 U3750 ( .A(a[20]), .ZN(n3109) );
  INV_X8 U3751 ( .A(b[3]), .ZN(n2506) );
  INV_X4 U3752 ( .A(a[24]), .ZN(n3589) );
  INV_X4 U3753 ( .A(n2785), .ZN(n3122) );
  INV_X4 U3754 ( .A(b[14]), .ZN(n2907) );
  NOR2_X4 U3755 ( .A1(n3010), .A2(n2907), .ZN(n2830) );
  MUX2_X2 U3756 ( .A(n1721), .B(n3208), .S(n94), .Z(n2480) );
  INV_X4 U3757 ( .A(a[19]), .ZN(n2407) );
  BUF_X4 U3758 ( .A(n2924), .Z(n2997) );
  OAI22_X2 U3760 ( .A1(n2997), .A2(n2415), .B1(n2414), .B2(n92), .ZN(n2418) );
  NOR2_X2 U3762 ( .A1(n2420), .A2(n2419), .ZN(n2508) );
  INV_X4 U3763 ( .A(a[21]), .ZN(n3217) );
  NOR2_X2 U3764 ( .A1(n2425), .A2(n602), .ZN(n2426) );
  INV_X4 U3766 ( .A(n97), .ZN(n2941) );
  NAND2_X2 U3768 ( .A1(n117), .A2(a[13]), .ZN(n2437) );
  NAND2_X1 U3769 ( .A1(n3329), .A2(n2407), .ZN(n2444) );
  NAND2_X2 U3770 ( .A1(n2450), .A2(n2449), .ZN(n2452) );
  NOR2_X2 U3771 ( .A1(n2454), .A2(n2455), .ZN(n2596) );
  INV_X4 U3772 ( .A(n2454), .ZN(n2457) );
  NOR2_X4 U3773 ( .A1(n2457), .A2(n2456), .ZN(n2597) );
  NAND2_X2 U3774 ( .A1(n2459), .A2(n2458), .ZN(n2461) );
  MUX2_X2 U3775 ( .A(n3310), .B(n3311), .S(a[22]), .Z(n2460) );
  NAND2_X2 U3776 ( .A1(n2461), .A2(n2460), .ZN(n2595) );
  MUX2_X2 U3777 ( .A(n1721), .B(n3208), .S(n96), .Z(n2478) );
  MUX2_X2 U3779 ( .A(n3203), .B(n1361), .S(n2941), .Z(n2467) );
  NAND2_X2 U3780 ( .A1(n2467), .A2(n2466), .ZN(n2468) );
  OAI21_X2 U3782 ( .B1(n2489), .B2(n2488), .A(n2487), .ZN(n2493) );
  MUX2_X2 U3783 ( .A(n1237), .B(n1381), .S(a[20]), .Z(n2494) );
  NAND2_X2 U3784 ( .A1(n2497), .A2(n2496), .ZN(n2588) );
  INV_X4 U3785 ( .A(a[13]), .ZN(n3202) );
  NAND2_X2 U3787 ( .A1(n2537), .A2(n2536), .ZN(n2540) );
  NAND2_X2 U3788 ( .A1(n2538), .A2(n3209), .ZN(n2539) );
  MUX2_X2 U3789 ( .A(n3311), .B(n3310), .S(n1554), .Z(n2548) );
  MUX2_X2 U3790 ( .A(n1303), .B(n3204), .S(n94), .Z(n2553) );
  INV_X4 U3792 ( .A(b[0]), .ZN(n3176) );
  NOR2_X2 U3794 ( .A1(n3303), .A2(a[23]), .ZN(n2558) );
  MUX2_X2 U3796 ( .A(n3203), .B(n3080), .S(n3109), .Z(n2574) );
  MUX2_X2 U3797 ( .A(n1303), .B(n3204), .S(a[19]), .Z(n2573) );
  NAND2_X2 U3798 ( .A1(n2574), .A2(n2573), .ZN(n2633) );
  NAND2_X2 U3799 ( .A1(n2578), .A2(n2577), .ZN(n2618) );
  MUX2_X2 U3800 ( .A(n3839), .B(n3113), .S(n3124), .Z(n2619) );
  XNOR2_X2 U3801 ( .A(n2618), .B(n2619), .ZN(n2579) );
  INV_X4 U3802 ( .A(n2581), .ZN(n2582) );
  AOI21_X2 U3803 ( .B1(n2583), .B2(n2251), .A(n2582), .ZN(n2647) );
  INV_X2 U3804 ( .A(n2585), .ZN(n2586) );
  MUX2_X2 U3805 ( .A(n3323), .B(n3329), .S(n2697), .Z(n2590) );
  INV_X2 U3806 ( .A(n2590), .ZN(n2592) );
  NOR2_X2 U3807 ( .A1(n2608), .A2(n2607), .ZN(n2612) );
  MUX2_X2 U3808 ( .A(n3839), .B(n3113), .S(a[17]), .Z(n2611) );
  INV_X4 U3809 ( .A(a[25]), .ZN(n2613) );
  AOI22_X2 U3810 ( .A1(n2622), .A2(n2621), .B1(n2620), .B2(n2619), .ZN(n2624)
         );
  NOR2_X2 U3811 ( .A1(n2625), .A2(n2624), .ZN(n2672) );
  INV_X4 U3812 ( .A(n2646), .ZN(n2644) );
  NOR2_X2 U3813 ( .A1(n2637), .A2(n2636), .ZN(n2666) );
  NAND2_X2 U3814 ( .A1(n2639), .A2(n2638), .ZN(n2667) );
  MUX2_X2 U3815 ( .A(n3203), .B(n84), .S(n3217), .Z(n2641) );
  NAND2_X2 U3817 ( .A1(n2641), .A2(n2640), .ZN(n2668) );
  XNOR2_X2 U3818 ( .A(n2666), .B(n2642), .ZN(n2645) );
  MUX2_X2 U3819 ( .A(n3323), .B(n3329), .S(n3589), .Z(n2658) );
  MUX2_X2 U3820 ( .A(n1237), .B(n1381), .S(a[23]), .Z(n2657) );
  MUX2_X2 U3822 ( .A(n3203), .B(n1361), .S(n2697), .Z(n2660) );
  MUX2_X2 U3823 ( .A(n1303), .B(n3204), .S(a[21]), .Z(n2659) );
  MUX2_X2 U3824 ( .A(a[25]), .B(b[7]), .S(n3132), .Z(n2662) );
  INV_X4 U3825 ( .A(n2760), .ZN(n2756) );
  MUX2_X2 U3826 ( .A(n1303), .B(n3204), .S(a[24]), .Z(n2680) );
  MUX2_X2 U3827 ( .A(n3839), .B(n3113), .S(a[21]), .Z(n2731) );
  XNOR2_X2 U3828 ( .A(n3595), .B(n2731), .ZN(n2685) );
  XNOR2_X2 U3829 ( .A(n2685), .B(n2684), .ZN(n2695) );
  MUX2_X2 U3830 ( .A(n3323), .B(n3329), .S(n2613), .Z(n2687) );
  NAND2_X2 U3832 ( .A1(n2687), .A2(n2686), .ZN(n2753) );
  MUX2_X2 U3833 ( .A(n2109), .B(n3208), .S(a[20]), .Z(n2715) );
  NOR2_X2 U3835 ( .A1(n2695), .A2(n2694), .ZN(n2730) );
  INV_X2 U3836 ( .A(n2730), .ZN(n2696) );
  NAND2_X2 U3837 ( .A1(n2695), .A2(n2694), .ZN(n2728) );
  NAND2_X2 U3838 ( .A1(n2696), .A2(n2728), .ZN(n2709) );
  MUX2_X2 U3839 ( .A(n3839), .B(n3113), .S(a[19]), .Z(n2700) );
  OAI21_X2 U3840 ( .B1(n2750), .B2(n2701), .A(n2751), .ZN(n2712) );
  MUX2_X2 U3841 ( .A(n2737), .B(n2736), .S(a[22]), .Z(n2703) );
  NOR2_X2 U3842 ( .A1(n2703), .A2(n2702), .ZN(n2707) );
  NAND2_X2 U3843 ( .A1(n2707), .A2(n2706), .ZN(n2710) );
  XOR2_X2 U3844 ( .A(n2709), .B(n2729), .Z(n3869) );
  XNOR2_X2 U3845 ( .A(n2713), .B(n2712), .ZN(n2727) );
  NOR2_X2 U3846 ( .A1(n2727), .A2(n2726), .ZN(n2745) );
  NOR2_X2 U3848 ( .A1(n3869), .A2(n3874), .ZN(n3682) );
  OAI22_X2 U3849 ( .A1(n2735), .A2(n2734), .B1(n2733), .B2(n2732), .ZN(n3582)
         );
  XNOR2_X2 U3850 ( .A(n3582), .B(n3583), .ZN(n2744) );
  MUX2_X2 U3851 ( .A(n2109), .B(n3208), .S(a[22]), .Z(n3593) );
  XNOR2_X2 U3853 ( .A(n2744), .B(n3581), .ZN(n3579) );
  NOR2_X2 U3854 ( .A1(n3580), .A2(n3579), .ZN(n3875) );
  NOR2_X2 U3855 ( .A1(n3682), .A2(n3875), .ZN(n2776) );
  INV_X1 U3856 ( .A(n2764), .ZN(n2755) );
  NOR2_X2 U3857 ( .A1(n1463), .A2(n2757), .ZN(n2761) );
  NOR2_X2 U3860 ( .A1(n2761), .A2(n2764), .ZN(n2762) );
  AOI21_X2 U3861 ( .B1(n2764), .B2(n1462), .A(n2762), .ZN(n2765) );
  BUF_X4 U3862 ( .A(n433), .Z(n2770) );
  NAND2_X2 U3863 ( .A1(n2776), .A2(n14), .ZN(n3617) );
  BUF_X4 U3864 ( .A(a[6]), .Z(n2906) );
  NAND2_X2 U3865 ( .A1(n2781), .A2(n2780), .ZN(n2791) );
  NAND2_X2 U3866 ( .A1(n3204), .A2(a[7]), .ZN(n2783) );
  INV_X4 U3867 ( .A(a[7]), .ZN(n3407) );
  NAND2_X2 U3868 ( .A1(n2783), .A2(n2782), .ZN(n2790) );
  NAND2_X2 U3869 ( .A1(n2785), .A2(b[4]), .ZN(n2802) );
  NAND2_X1 U3870 ( .A1(n3203), .A2(a[7]), .ZN(n2792) );
  NOR2_X2 U3871 ( .A1(n2145), .A2(n3498), .ZN(n2803) );
  NOR2_X2 U3874 ( .A1(n2803), .A2(n2800), .ZN(n2801) );
  NOR2_X2 U3875 ( .A1(n2858), .A2(n2814), .ZN(n2861) );
  NOR2_X2 U3876 ( .A1(n2813), .A2(n2858), .ZN(n2811) );
  NOR2_X2 U3877 ( .A1(n2861), .A2(n2811), .ZN(n2818) );
  BUF_X4 U3878 ( .A(a[5]), .Z(n3389) );
  INV_X4 U3879 ( .A(n2819), .ZN(n3392) );
  BUF_X4 U3880 ( .A(b[1]), .Z(n2983) );
  NAND2_X1 U3881 ( .A1(n3118), .A2(n3003), .ZN(n2831) );
  NOR2_X2 U3883 ( .A1(n2833), .A2(n2832), .ZN(n2834) );
  NOR2_X2 U3884 ( .A1(n2926), .A2(n2927), .ZN(n2844) );
  NOR2_X2 U3885 ( .A1(n2841), .A2(n602), .ZN(n2842) );
  NAND2_X2 U3886 ( .A1(n1721), .A2(n2355), .ZN(n2848) );
  NAND2_X2 U3887 ( .A1(n2863), .A2(n2862), .ZN(n2864) );
  BUF_X4 U3888 ( .A(a[6]), .Z(n3468) );
  MUX2_X2 U3889 ( .A(n1303), .B(n3204), .S(n1652), .Z(n2866) );
  NAND2_X2 U3890 ( .A1(n2867), .A2(n2866), .ZN(n2868) );
  NAND2_X2 U3891 ( .A1(n249), .A2(a[3]), .ZN(n2871) );
  AOI21_X2 U3893 ( .B1(n2904), .B2(n2905), .A(n1685), .ZN(n2936) );
  INV_X4 U3894 ( .A(a[0]), .ZN(n2998) );
  INV_X4 U3895 ( .A(n2998), .ZN(n3515) );
  NAND2_X2 U3896 ( .A1(n2896), .A2(n2895), .ZN(n2990) );
  NAND2_X2 U3897 ( .A1(n3119), .A2(n99), .ZN(n2898) );
  NAND2_X2 U3898 ( .A1(n2898), .A2(n2897), .ZN(n2900) );
  OAI22_X2 U3900 ( .A1(n2909), .A2(n2997), .B1(n92), .B2(n2908), .ZN(n2912) );
  MUX2_X2 U3902 ( .A(n3119), .B(n3120), .S(n56), .Z(n2957) );
  NOR2_X2 U3904 ( .A1(n3323), .A2(n3202), .ZN(n2938) );
  MUX2_X2 U3906 ( .A(n3454), .B(n3455), .S(n2400), .Z(n2942) );
  MUX2_X2 U3907 ( .A(n3311), .B(n3310), .S(n2438), .Z(n3194) );
  INV_X4 U3908 ( .A(n2190), .ZN(n2959) );
  BUF_X4 U3909 ( .A(n2968), .Z(n2969) );
  AOI21_X2 U3910 ( .B1(n3177), .B2(n916), .A(n2997), .ZN(n3000) );
  INV_X4 U3911 ( .A(n2998), .ZN(n3538) );
  MUX2_X2 U3912 ( .A(n988), .B(n2315), .S(n1221), .Z(n3006) );
  NAND3_X2 U3913 ( .A1(n3011), .A2(n92), .A3(n4149), .ZN(n3057) );
  MUX2_X2 U3914 ( .A(n1303), .B(n3204), .S(n2356), .Z(n3028) );
  AOI22_X2 U3915 ( .A1(n3019), .A2(n34), .B1(n77), .B2(n3018), .ZN(n3090) );
  NAND2_X2 U3916 ( .A1(n3029), .A2(n3028), .ZN(n3031) );
  MUX2_X2 U3917 ( .A(n3513), .B(n1407), .S(a[12]), .Z(n3036) );
  INV_X2 U3918 ( .A(n3301), .ZN(n3078) );
  OAI21_X2 U3919 ( .B1(n1314), .B2(n3362), .A(n3361), .ZN(n3372) );
  INV_X4 U3920 ( .A(n3094), .ZN(n3101) );
  BUF_X4 U3921 ( .A(n3097), .Z(n3098) );
  XNOR2_X2 U3923 ( .A(n97), .B(n3122), .ZN(n3123) );
  NAND2_X2 U3924 ( .A1(n3155), .A2(n1238), .ZN(n3138) );
  NAND2_X2 U3925 ( .A1(n3145), .A2(n3148), .ZN(n3151) );
  NOR3_X2 U3927 ( .A1(n3163), .A2(n2230), .A3(n1788), .ZN(n3167) );
  NOR2_X2 U3928 ( .A1(n3163), .A2(n2230), .ZN(n3166) );
  OAI22_X2 U3929 ( .A1(n3167), .A2(n454), .B1(n3166), .B2(n3165), .ZN(n3169)
         );
  MUX2_X2 U3930 ( .A(n3455), .B(n3454), .S(n97), .Z(n3201) );
  MUX2_X2 U3931 ( .A(n2830), .B(n3208), .S(n56), .Z(n3216) );
  OAI22_X2 U3932 ( .A1(n3212), .A2(n3211), .B1(n3306), .B2(n3210), .ZN(n3215)
         );
  NAND2_X2 U3934 ( .A1(n3295), .A2(n3249), .ZN(n3225) );
  OAI21_X2 U3935 ( .B1(n414), .B2(n3223), .A(n3222), .ZN(n3293) );
  NOR2_X2 U3937 ( .A1(n56), .A2(n3303), .ZN(n3304) );
  NOR2_X2 U3938 ( .A1(n3307), .A2(n3306), .ZN(n3308) );
  MUX2_X2 U3939 ( .A(n3311), .B(n3310), .S(n3534), .Z(n3384) );
  NOR2_X2 U3941 ( .A1(n3320), .A2(n3319), .ZN(n3347) );
  MUX2_X2 U3942 ( .A(n3323), .B(n3329), .S(n2045), .Z(n3325) );
  MUX2_X2 U3943 ( .A(n1237), .B(n1381), .S(n3538), .Z(n3324) );
  NAND2_X2 U3944 ( .A1(n3325), .A2(n3324), .ZN(n3388) );
  MUX2_X2 U3945 ( .A(n3513), .B(n1407), .S(a[9]), .Z(n3327) );
  XNOR2_X2 U3946 ( .A(n3344), .B(n3343), .ZN(n3345) );
  INV_X4 U3947 ( .A(n3372), .ZN(n3373) );
  MUX2_X2 U3948 ( .A(n1262), .B(n3454), .S(n2356), .Z(n3405) );
  NOR2_X2 U3949 ( .A1(n3406), .A2(n3405), .ZN(n3464) );
  INV_X4 U3950 ( .A(n3463), .ZN(n3423) );
  NAND2_X2 U3951 ( .A1(n3411), .A2(n3410), .ZN(n3412) );
  NOR2_X2 U3952 ( .A1(n3415), .A2(n3414), .ZN(n3422) );
  NAND2_X2 U3953 ( .A1(n3426), .A2(n3425), .ZN(n3429) );
  MUX2_X2 U3954 ( .A(n1209), .B(n1863), .S(n99), .Z(n3432) );
  MUX2_X2 U3955 ( .A(n3455), .B(n3454), .S(a[1]), .Z(n3456) );
  NOR2_X2 U3956 ( .A1(n3457), .A2(n3456), .ZN(n3466) );
  MUX2_X2 U3957 ( .A(n1266), .B(n3522), .S(n3534), .Z(n3461) );
  AND3_X1 U3958 ( .A1(n3480), .A2(n3482), .A3(n3487), .ZN(n3481) );
  NAND2_X2 U3959 ( .A1(n3474), .A2(n3473), .ZN(n3544) );
  MUX2_X2 U3960 ( .A(n3513), .B(n3512), .S(n1221), .Z(n3478) );
  NAND2_X2 U3961 ( .A1(n3478), .A2(n3477), .ZN(n3537) );
  NAND2_X2 U3962 ( .A1(n3544), .A2(n3537), .ZN(n3545) );
  INV_X2 U3963 ( .A(n3487), .ZN(n3490) );
  AOI22_X2 U3964 ( .A1(n3490), .A2(n3489), .B1(n3488), .B2(n3487), .ZN(n3769)
         );
  NOR2_X2 U3965 ( .A1(n1672), .A2(n1666), .ZN(n3491) );
  NOR2_X1 U3966 ( .A1(n3532), .A2(n3495), .ZN(n3497) );
  OAI22_X2 U3968 ( .A1(n3520), .A2(n3519), .B1(n1649), .B2(n3518), .ZN(n3523)
         );
  NAND3_X2 U3969 ( .A1(n3523), .A2(n3522), .A3(n3521), .ZN(n3524) );
  NOR2_X1 U3970 ( .A1(n3528), .A2(n3527), .ZN(n3530) );
  INV_X1 U3972 ( .A(n3530), .ZN(n3531) );
  AOI22_X2 U3973 ( .A1(n3533), .A2(n3532), .B1(n1147), .B2(n3531), .ZN(n3541)
         );
  XNOR2_X2 U3974 ( .A(n3550), .B(n3544), .ZN(n3540) );
  INV_X1 U3977 ( .A(n3545), .ZN(n3546) );
  AOI21_X2 U3978 ( .B1(n3548), .B2(n3547), .A(n3546), .ZN(n3554) );
  OAI22_X2 U3979 ( .A1(n3554), .A2(n3553), .B1(n3552), .B2(n3551), .ZN(n3762)
         );
  INV_X4 U3980 ( .A(n3720), .ZN(n3710) );
  NOR2_X4 U3981 ( .A1(n3909), .A2(n3910), .ZN(n4010) );
  NAND2_X2 U3982 ( .A1(n3869), .A2(n3874), .ZN(n3683) );
  INV_X2 U3983 ( .A(n3875), .ZN(n3868) );
  NAND2_X2 U3986 ( .A1(n3664), .A2(n3866), .ZN(n3619) );
  MUX2_X2 U3987 ( .A(n2109), .B(n3208), .S(a[23]), .Z(n3645) );
  INV_X4 U3988 ( .A(n4021), .ZN(n3730) );
  NOR2_X4 U3990 ( .A1(n3714), .A2(n3709), .ZN(n3678) );
  NAND2_X2 U3991 ( .A1(n3678), .A2(n3616), .ZN(n3635) );
  NAND2_X2 U3992 ( .A1(n3678), .A2(n3628), .ZN(n3629) );
  OAI22_X2 U3993 ( .A1(n3924), .A2(n3629), .B1(n3678), .B2(n3628), .ZN(n3630)
         );
  AOI21_X2 U3994 ( .B1(n3631), .B2(n1804), .A(n3630), .ZN(n3632) );
  NOR2_X1 U3995 ( .A1(n3639), .A2(n3646), .ZN(n3642) );
  INV_X1 U3998 ( .A(n3645), .ZN(n3649) );
  NOR2_X1 U3999 ( .A1(n3650), .A2(n3649), .ZN(n3653) );
  INV_X1 U4000 ( .A(n3651), .ZN(n3652) );
  NOR2_X2 U4001 ( .A1(n3656), .A2(n2388), .ZN(n3657) );
  NAND4_X1 U4002 ( .A1(n3683), .A2(n3711), .A3(n1586), .A4(n3663), .ZN(n3660)
         );
  INV_X1 U4003 ( .A(n3668), .ZN(n3665) );
  INV_X2 U4004 ( .A(n3675), .ZN(n3687) );
  NAND2_X2 U4005 ( .A1(n3866), .A2(n3868), .ZN(n3680) );
  NAND3_X2 U4006 ( .A1(n3687), .A2(n3683), .A3(n3680), .ZN(n3679) );
  NAND2_X2 U4007 ( .A1(n3678), .A2(n3676), .ZN(n3693) );
  INV_X4 U4008 ( .A(n14), .ZN(n3919) );
  NOR3_X2 U4009 ( .A1(n3919), .A2(n3682), .A3(n3680), .ZN(n3685) );
  NOR2_X2 U4011 ( .A1(n3678), .A2(n3677), .ZN(n3692) );
  NOR2_X2 U4012 ( .A1(n3679), .A2(n3710), .ZN(n3691) );
  INV_X2 U4013 ( .A(n3680), .ZN(n3681) );
  NOR2_X1 U4015 ( .A1(n3917), .A2(n3919), .ZN(n3688) );
  OAI22_X2 U4016 ( .A1(n3689), .A2(n3688), .B1(n3687), .B2(n3686), .ZN(n3690)
         );
  AOI21_X2 U4017 ( .B1(n1804), .B2(n3695), .A(n3694), .ZN(n3697) );
  NAND2_X2 U4018 ( .A1(n3698), .A2(n3722), .ZN(n3701) );
  AOI21_X2 U4019 ( .B1(n3710), .B2(n3709), .A(n3708), .ZN(n3718) );
  OAI211_X1 U4020 ( .C1(n3725), .C2(n3729), .A(n3724), .B(n3723), .ZN(n3726)
         );
  NOR2_X2 U4021 ( .A1(n3727), .A2(n3726), .ZN(n3733) );
  NAND2_X2 U4023 ( .A1(n3741), .A2(n3740), .ZN(n3744) );
  NAND2_X2 U4024 ( .A1(n3744), .A2(n3743), .ZN(\d[25] ) );
  NOR2_X2 U4025 ( .A1(n3748), .A2(n1380), .ZN(n3754) );
  INV_X4 U4026 ( .A(n3749), .ZN(n3820) );
  NOR2_X2 U4027 ( .A1(n3820), .A2(n3750), .ZN(n3751) );
  NAND2_X2 U4028 ( .A1(n3751), .A2(n3833), .ZN(n3752) );
  BUF_X4 U4029 ( .A(n3829), .Z(n3904) );
  INV_X4 U4030 ( .A(n3904), .ZN(n3794) );
  OAI21_X2 U4031 ( .B1(n3890), .B2(n3887), .A(n3755), .ZN(n3977) );
  BUF_X4 U4032 ( .A(n3776), .Z(n3784) );
  XNOR2_X2 U4033 ( .A(n3790), .B(n3789), .ZN(\d[13]_BAR ) );
  NAND2_X2 U4035 ( .A1(n3796), .A2(n3795), .ZN(\d[16]_BAR ) );
  XNOR2_X2 U4036 ( .A(n3802), .B(n3801), .ZN(\d[14]_BAR ) );
  OAI22_X2 U4037 ( .A1(n3819), .A2(n3818), .B1(n3817), .B2(n3816), .ZN(n3822)
         );
  NAND2_X2 U4040 ( .A1(n3873), .A2(n3880), .ZN(n3870) );
  BUF_X4 U4041 ( .A(n3883), .Z(n3884) );
  NAND2_X2 U4043 ( .A1(n3886), .A2(n3887), .ZN(n3901) );
  OAI211_X1 U4044 ( .C1(n3901), .C2(n891), .A(n3900), .B(n3899), .ZN(n3902) );
  NOR2_X2 U4045 ( .A1(n3903), .A2(n3902), .ZN(\d[21]_BAR ) );
  MUX2_X2 U4046 ( .A(n3961), .B(n1787), .S(n3912), .Z(n3913) );
  INV_X4 U4047 ( .A(n3929), .ZN(n3927) );
  OAI21_X2 U4048 ( .B1(n3924), .B2(n3923), .A(n3922), .ZN(n3925) );
  AOI21_X2 U4049 ( .B1(n3927), .B2(n3926), .A(n3925), .ZN(n3931) );
  NOR2_X2 U4050 ( .A1(n3934), .A2(n1482), .ZN(n3944) );
  NAND2_X2 U4051 ( .A1(n3935), .A2(n4015), .ZN(n3943) );
  NAND2_X2 U4053 ( .A1(n3952), .A2(n3951), .ZN(\d[24]_BAR ) );
  NAND4_X1 U4054 ( .A1(n3971), .A2(n3970), .A3(n4010), .A4(n3969), .ZN(n3972)
         );
  NAND3_X2 U4055 ( .A1(n3974), .A2(n3972), .A3(n3973), .ZN(n3975) );
  AOI21_X2 U4056 ( .B1(n3977), .B2(n3976), .A(n3975), .ZN(n3980) );
  NOR2_X2 U4057 ( .A1(n3995), .A2(n4018), .ZN(n3997) );
  NAND3_X2 U4058 ( .A1(n4002), .A2(n4001), .A3(n4000), .ZN(\d[30]_BAR ) );
  OAI22_X2 U4059 ( .A1(n4022), .A2(n4015), .B1(n4020), .B2(n4021), .ZN(n4027)
         );
  NAND2_X2 U2306 ( .A1(n831), .A2(n2045), .ZN(n3426) );
  NAND2_X4 U994 ( .A1(n252), .A2(n251), .ZN(n572) );
  NAND2_X4 U995 ( .A1(b[11]), .A2(b[12]), .ZN(n251) );
  NOR2_X4 U866 ( .A1(n2005), .A2(n220), .ZN(n1912) );
  NAND2_X4 U2275 ( .A1(n3244), .A2(n3245), .ZN(n3243) );
  INV_X2 U934 ( .A(n2812), .ZN(n233) );
  NAND2_X2 U26 ( .A1(n97), .A2(n1478), .ZN(n1338) );
  NAND2_X2 U2865 ( .A1(n1766), .A2(n3109), .ZN(n2224) );
  INV_X2 U2856 ( .A(n3303), .ZN(n1859) );
  NAND2_X2 U2741 ( .A1(n1210), .A2(n1211), .ZN(n1213) );
  INV_X1 U200 ( .A(n3963), .ZN(n520) );
  NAND2_X2 U2740 ( .A1(n3134), .A2(n2187), .ZN(n1212) );
  NAND2_X4 U7 ( .A1(n1559), .A2(n1560), .ZN(n1562) );
  NOR2_X4 U483 ( .A1(n73), .A2(n1557), .ZN(n109) );
  NAND2_X4 U1173 ( .A1(n349), .A2(n2655), .ZN(n2772) );
  NAND2_X2 U3012 ( .A1(n3376), .A2(n3375), .ZN(n3379) );
  NAND2_X2 U306 ( .A1(n1254), .A2(n2756), .ZN(n1256) );
  INV_X4 U254 ( .A(n3709), .ZN(n3698) );
  NAND2_X2 U307 ( .A1(n741), .A2(n740), .ZN(n391) );
  INV_X2 U2007 ( .A(n2559), .ZN(n617) );
  NAND2_X4 U1234 ( .A1(n3258), .A2(n3257), .ZN(n3282) );
  NAND2_X4 U1178 ( .A1(n352), .A2(n351), .ZN(n2974) );
  NAND2_X2 U501 ( .A1(n97), .A2(n111), .ZN(n2071) );
  INV_X4 U2812 ( .A(n1209), .ZN(n1266) );
  NOR2_X2 U2704 ( .A1(n1197), .A2(n3062), .ZN(n1196) );
  INV_X4 U2411 ( .A(n244), .ZN(n2816) );
  INV_X4 U1040 ( .A(n3177), .ZN(n3008) );
  INV_X4 U337 ( .A(n2018), .ZN(n1441) );
  AND2_X2 U115 ( .A1(n2982), .A2(a[14]), .ZN(n15) );
  NAND3_X2 U2588 ( .A1(n1337), .A2(n57), .A3(n55), .ZN(n1092) );
  NAND2_X1 U1471 ( .A1(n1149), .A2(n3529), .ZN(n1148) );
  NAND2_X2 U1497 ( .A1(n3526), .A2(n3524), .ZN(n1674) );
  INV_X4 U2281 ( .A(n892), .ZN(n810) );
  NAND2_X2 U167 ( .A1(n47), .A2(n44), .ZN(n2608) );
  INV_X2 U2317 ( .A(n2655), .ZN(n848) );
  AOI22_X2 U3291 ( .A1(n3034), .A2(a[8]), .B1(n249), .B2(a[7]), .ZN(n2144) );
  NOR2_X4 U925 ( .A1(b[11]), .A2(b[12]), .ZN(n253) );
  NAND2_X1 U3926 ( .A1(n3148), .A2(n3147), .ZN(n3149) );
  INV_X2 U191 ( .A(n3154), .ZN(n3144) );
  XNOR2_X1 U4014 ( .A(n3683), .B(n3681), .ZN(n3689) );
  NAND2_X2 U3791 ( .A1(n2736), .A2(a[12]), .ZN(n2555) );
  NAND2_X4 U605 ( .A1(n2423), .A2(b[8]), .ZN(n156) );
  NAND2_X2 U245 ( .A1(n3848), .A2(n3668), .ZN(n3661) );
  INV_X4 U3595 ( .A(a[15]), .ZN(n2079) );
  AOI22_X2 U1565 ( .A1(n3119), .A2(n2258), .B1(n3120), .B2(a[11]), .ZN(n1117)
         );
  INV_X4 U2754 ( .A(n216), .ZN(n3961) );
  NOR2_X4 U724 ( .A1(n1113), .A2(n2006), .ZN(n2005) );
  NOR2_X4 U2903 ( .A1(n2596), .A2(n2597), .ZN(n2462) );
  NAND2_X1 U1390 ( .A1(n249), .A2(a[10]), .ZN(n3179) );
  NAND2_X2 U1636 ( .A1(n2581), .A2(n2583), .ZN(n1136) );
  AOI22_X2 U155 ( .A1(n3881), .A2(n147), .B1(n3879), .B2(n3880), .ZN(n3882) );
  NAND2_X2 U1587 ( .A1(n2481), .A2(n2158), .ZN(n1430) );
  NAND2_X2 U2885 ( .A1(n2868), .A2(n2869), .ZN(n2893) );
  NAND2_X2 U681 ( .A1(n519), .A2(n76), .ZN(n1460) );
  OAI22_X2 U3669 ( .A1(n2290), .A2(n1471), .B1(n3720), .B2(n4079), .ZN(n3562)
         );
  INV_X4 U3088 ( .A(n2556), .ZN(n2198) );
  NAND2_X2 U1657 ( .A1(n955), .A2(n710), .ZN(n629) );
  NAND2_X2 U3511 ( .A1(n1863), .A2(n3202), .ZN(n1920) );
  NAND2_X4 U543 ( .A1(n931), .A2(n3933), .ZN(n2000) );
  NOR2_X2 U1380 ( .A1(n3699), .A2(n3612), .ZN(n2679) );
  INV_X4 U2456 ( .A(n2948), .ZN(n972) );
  NAND2_X4 U575 ( .A1(n3563), .A2(n3562), .ZN(n147) );
  INV_X4 U2069 ( .A(n1926), .ZN(n621) );
  INV_X2 U281 ( .A(n2584), .ZN(n1267) );
  INV_X2 U428 ( .A(n2982), .ZN(n91) );
  NOR2_X2 U3736 ( .A1(n3915), .A2(n3916), .ZN(n3926) );
  NAND2_X2 U3208 ( .A1(n2220), .A2(n2789), .ZN(n2215) );
  NAND3_X2 U1658 ( .A1(n2048), .A2(n803), .A3(n2218), .ZN(n627) );
  INV_X4 U2259 ( .A(n2116), .ZN(n790) );
  INV_X4 U2065 ( .A(n1569), .ZN(n618) );
  NAND2_X4 U1973 ( .A1(n560), .A2(n1057), .ZN(n2789) );
  NAND2_X2 U1953 ( .A1(n1180), .A2(n2513), .ZN(n545) );
  INV_X2 U25 ( .A(n2051), .ZN(n1393) );
  INV_X4 U2112 ( .A(n1299), .ZN(n653) );
  INV_X2 U3901 ( .A(n2916), .ZN(n2918) );
  NAND2_X1 U3971 ( .A1(n3529), .A2(n3530), .ZN(n3533) );
  AOI21_X2 U1756 ( .B1(n3524), .B2(n3525), .A(n74), .ZN(n1673) );
  NOR2_X4 U2623 ( .A1(n2115), .A2(n1123), .ZN(n1869) );
  NAND2_X4 U902 ( .A1(n791), .A2(n790), .ZN(n2115) );
  INV_X2 U2152 ( .A(n710), .ZN(n954) );
  NOR3_X1 U3136 ( .A1(n3067), .A2(n2506), .A3(a[15]), .ZN(n2826) );
  NAND2_X2 U159 ( .A1(n3068), .A2(n1478), .ZN(n33) );
  INV_X4 U3496 ( .A(n3066), .ZN(n3067) );
  INV_X2 U169 ( .A(a[23]), .ZN(n45) );
  INV_X4 U433 ( .A(n2442), .ZN(n97) );
  INV_X4 U1871 ( .A(n481), .ZN(n3453) );
  NAND2_X2 U809 ( .A1(n3034), .A2(n1837), .ZN(n2022) );
  INV_X4 U2565 ( .A(n3454), .ZN(n3472) );
  NOR2_X2 U2878 ( .A1(n2550), .A2(n2549), .ZN(n2552) );
  NOR2_X2 U3303 ( .A1(n1954), .A2(n3201), .ZN(n3239) );
  NAND2_X2 U819 ( .A1(n207), .A2(n2996), .ZN(n1729) );
  NOR2_X2 U3218 ( .A1(n2452), .A2(n2451), .ZN(n2454) );
  NAND2_X2 U1898 ( .A1(n1863), .A2(n2228), .ZN(n503) );
  NAND2_X2 U3338 ( .A1(n2720), .A2(n2719), .ZN(n2764) );
  NOR2_X2 U2815 ( .A1(n3006), .A2(n3005), .ZN(n3062) );
  NAND2_X1 U3661 ( .A1(n2254), .A2(n465), .ZN(n2464) );
  NAND2_X2 U183 ( .A1(n367), .A2(n263), .ZN(n366) );
  NOR2_X2 U1205 ( .A1(n371), .A2(n2541), .ZN(n3291) );
  NAND2_X2 U9 ( .A1(n3170), .A2(n2317), .ZN(n1038) );
  NOR2_X2 U3122 ( .A1(n2674), .A2(n2672), .ZN(n2630) );
  NAND2_X2 U1864 ( .A1(n477), .A2(n478), .ZN(n2601) );
  NAND2_X2 U864 ( .A1(n1563), .A2(n1564), .ZN(n218) );
  INV_X4 U1800 ( .A(a[10]), .ZN(n2228) );
  NAND2_X2 U3 ( .A1(n1412), .A2(n1413), .ZN(n3578) );
  NOR2_X2 U5 ( .A1(n491), .A2(n492), .ZN(n415) );
  INV_X4 U10 ( .A(n4099), .ZN(n241) );
  NAND2_X2 U12 ( .A1(n1337), .A2(n54), .ZN(n1339) );
  NOR2_X2 U13 ( .A1(n3303), .A2(a[19]), .ZN(n2923) );
  AND2_X1 U14 ( .A1(n2315), .A2(n88), .ZN(n458) );
  NOR2_X1 U17 ( .A1(n1303), .A2(n55), .ZN(n327) );
  NAND2_X1 U20 ( .A1(n881), .A2(n880), .ZN(n197) );
  OR2_X1 U21 ( .A1(n3589), .A2(n3498), .ZN(n456) );
  OR2_X1 U22 ( .A1(n85), .A2(n97), .ZN(n16) );
  NAND2_X1 U31 ( .A1(n2917), .A2(n2916), .ZN(n777) );
  NAND2_X2 U38 ( .A1(n4127), .A2(n1879), .ZN(n1629) );
  NAND2_X1 U39 ( .A1(n2962), .A2(n18), .ZN(n3161) );
  NAND2_X1 U41 ( .A1(n4045), .A2(a[12]), .ZN(n795) );
  NAND2_X1 U42 ( .A1(n2312), .A2(n2311), .ZN(n2433) );
  NAND2_X1 U48 ( .A1(a[24]), .A2(n3453), .ZN(n173) );
  NAND3_X1 U50 ( .A1(n632), .A2(n2131), .A3(n631), .ZN(n344) );
  NAND2_X1 U53 ( .A1(n4036), .A2(n859), .ZN(n858) );
  NAND2_X2 U54 ( .A1(n2552), .A2(n2551), .ZN(n272) );
  NAND2_X1 U55 ( .A1(n2736), .A2(a[20]), .ZN(n354) );
  NAND2_X1 U56 ( .A1(n2514), .A2(n2518), .ZN(n132) );
  INV_X1 U57 ( .A(n1211), .ZN(n2187) );
  INV_X1 U63 ( .A(n1116), .ZN(n1353) );
  MUX2_X1 U64 ( .A(n3513), .B(n3512), .S(a[3]), .Z(n3504) );
  INV_X4 U66 ( .A(n3176), .ZN(n2982) );
  MUX2_X1 U69 ( .A(n241), .B(n117), .S(n3124), .Z(n2496) );
  OR2_X1 U71 ( .A1(n733), .A2(n2478), .ZN(n465) );
  MUX2_X1 U76 ( .A(n86), .B(n2058), .S(n2697), .Z(n2607) );
  NAND2_X1 U80 ( .A1(n340), .A2(n344), .ZN(n343) );
  INV_X2 U81 ( .A(n2533), .ZN(n1375) );
  INV_X2 U91 ( .A(n1085), .ZN(n1514) );
  INV_X1 U93 ( .A(n3053), .ZN(n1422) );
  NOR2_X1 U94 ( .A1(n2429), .A2(n2428), .ZN(n2486) );
  NAND2_X1 U111 ( .A1(n2468), .A2(n2469), .ZN(n2474) );
  INV_X2 U116 ( .A(n1810), .ZN(n1563) );
  INV_X1 U117 ( .A(n3258), .ZN(n2330) );
  NAND2_X1 U122 ( .A1(n1377), .A2(n95), .ZN(n703) );
  INV_X1 U123 ( .A(n3332), .ZN(n2366) );
  NAND2_X2 U125 ( .A1(n1138), .A2(n2464), .ZN(n2581) );
  MUX2_X1 U134 ( .A(n2980), .B(n2022), .S(a[19]), .Z(n2639) );
  AOI21_X1 U137 ( .B1(n2967), .B2(n2969), .A(n2972), .ZN(n4197) );
  MUX2_X1 U138 ( .A(n1237), .B(n1381), .S(a[24]), .Z(n2686) );
  NAND2_X1 U139 ( .A1(n762), .A2(n2253), .ZN(n1872) );
  NAND2_X1 U140 ( .A1(n1766), .A2(n3407), .ZN(n1033) );
  MUX2_X1 U147 ( .A(n87), .B(n1121), .S(n1221), .Z(n3391) );
  NOR2_X2 U154 ( .A1(n1831), .A2(n3044), .ZN(n3022) );
  MUX2_X1 U157 ( .A(n2654), .B(n2296), .S(n3217), .Z(n2702) );
  INV_X1 U165 ( .A(n3232), .ZN(n4082) );
  OR2_X1 U179 ( .A1(n333), .A2(n1005), .ZN(n52) );
  OAI22_X1 U187 ( .A1(n2693), .A2(n2715), .B1(n2753), .B2(n2714), .ZN(n2694)
         );
  NAND2_X2 U211 ( .A1(n1740), .A2(n1741), .ZN(n1299) );
  BUF_X1 U246 ( .A(n3746), .Z(n4186) );
  NAND2_X1 U255 ( .A1(n3036), .A2(n3035), .ZN(n3343) );
  NAND2_X2 U264 ( .A1(n940), .A2(n2500), .ZN(n2603) );
  NAND2_X2 U273 ( .A1(n1003), .A2(n52), .ZN(n3095) );
  INV_X2 U275 ( .A(n1912), .ZN(n1528) );
  INV_X2 U284 ( .A(n1383), .ZN(n67) );
  INV_X1 U290 ( .A(n2653), .ZN(n893) );
  AOI22_X1 U294 ( .A1(n2606), .A2(n1156), .B1(n1155), .B2(n2603), .ZN(n1604)
         );
  NAND2_X2 U310 ( .A1(n763), .A2(n1604), .ZN(n4019) );
  NAND2_X2 U318 ( .A1(n1639), .A2(n4008), .ZN(n1617) );
  INV_X1 U324 ( .A(n3934), .ZN(n3939) );
  INV_X1 U326 ( .A(n2320), .ZN(n3804) );
  INV_X1 U333 ( .A(n61), .ZN(n2061) );
  NAND2_X2 U334 ( .A1(n1921), .A2(n3438), .ZN(n3781) );
  NOR2_X1 U358 ( .A1(n3905), .A2(n298), .ZN(n293) );
  XNOR2_X1 U372 ( .A(n3822), .B(n3821), .ZN(\d[15]_BAR ) );
  AND2_X1 U379 ( .A1(n3920), .A2(n3854), .ZN(n4031) );
  OR2_X1 U398 ( .A1(n2883), .A2(n2983), .ZN(n4033) );
  OR2_X1 U400 ( .A1(n3328), .A2(n93), .ZN(n4034) );
  NAND2_X1 U401 ( .A1(n2882), .A2(n3067), .ZN(n4035) );
  OR2_X1 U404 ( .A1(n3455), .A2(n56), .ZN(n4036) );
  OR2_X1 U405 ( .A1(n3200), .A2(n56), .ZN(n4037) );
  OR2_X1 U409 ( .A1(n4075), .A2(n3407), .ZN(n4038) );
  AND3_X1 U413 ( .A1(n1487), .A2(n1818), .A3(n3407), .ZN(n4039) );
  OR2_X2 U417 ( .A1(n2299), .A2(a[11]), .ZN(n4040) );
  OR2_X1 U419 ( .A1(n3200), .A2(a[11]), .ZN(n4041) );
  OR2_X1 U420 ( .A1(n3208), .A2(n2258), .ZN(n4042) );
  AND2_X1 U426 ( .A1(a[3]), .A2(n2924), .ZN(n4044) );
  INV_X2 U430 ( .A(a[1]), .ZN(n2045) );
  OAI21_X1 U434 ( .B1(n2845), .B2(n710), .A(n2013), .ZN(n2934) );
  INV_X1 U454 ( .A(n1311), .ZN(n3955) );
  AND2_X4 U456 ( .A1(n2741), .A2(n2742), .ZN(n4045) );
  AND2_X1 U459 ( .A1(n3003), .A2(n3413), .ZN(n4046) );
  AND2_X2 U461 ( .A1(n1995), .A2(n1992), .ZN(n4047) );
  OR2_X1 U467 ( .A1(a[17]), .A2(n1928), .ZN(n4049) );
  OR2_X1 U475 ( .A1(n2506), .A2(a[24]), .ZN(n4051) );
  AND2_X1 U477 ( .A1(n1766), .A2(n3589), .ZN(n4052) );
  OR2_X1 U478 ( .A1(n2980), .A2(a[14]), .ZN(n4053) );
  AND2_X2 U479 ( .A1(n2220), .A2(n2789), .ZN(n4054) );
  OR2_X1 U490 ( .A1(n602), .A2(n467), .ZN(n4055) );
  OR2_X1 U494 ( .A1(n3455), .A2(n98), .ZN(n4056) );
  OR2_X1 U506 ( .A1(n3008), .A2(a[12]), .ZN(n4057) );
  OR2_X1 U507 ( .A1(n3200), .A2(a[12]), .ZN(n4058) );
  OR2_X1 U518 ( .A1(a[23]), .A2(n3455), .ZN(n4059) );
  AND2_X1 U522 ( .A1(n3809), .A2(n2320), .ZN(n4060) );
  AND2_X1 U531 ( .A1(n313), .A2(n3515), .ZN(n4063) );
  INV_X4 U532 ( .A(n2400), .ZN(n3124) );
  INV_X2 U533 ( .A(a[8]), .ZN(n3413) );
  BUF_X1 U535 ( .A(n3287), .Z(n1631) );
  AND2_X2 U536 ( .A1(n872), .A2(n2812), .ZN(n4064) );
  BUF_X2 U541 ( .A(n1928), .Z(n3522) );
  INV_X2 U558 ( .A(n2881), .ZN(n1326) );
  INV_X1 U577 ( .A(n2580), .ZN(n2251) );
  AOI21_X1 U579 ( .B1(n2474), .B2(n2475), .A(n2472), .ZN(n2580) );
  AND2_X2 U580 ( .A1(n1045), .A2(n1162), .ZN(n4065) );
  INV_X2 U587 ( .A(a[12]), .ZN(n3016) );
  INV_X1 U591 ( .A(n414), .ZN(n3220) );
  INV_X2 U592 ( .A(a[3]), .ZN(n2026) );
  OR2_X1 U598 ( .A1(n1507), .A2(n3085), .ZN(n4066) );
  OR3_X1 U599 ( .A1(n1272), .A2(n70), .A3(n2368), .ZN(n4067) );
  OR2_X1 U600 ( .A1(n3371), .A2(n2088), .ZN(n4068) );
  INV_X2 U607 ( .A(n1840), .ZN(n2935) );
  OR2_X2 U608 ( .A1(n2309), .A2(n2501), .ZN(n4069) );
  AND2_X1 U609 ( .A1(n3998), .A2(n4010), .ZN(n4070) );
  AND2_X2 U622 ( .A1(n133), .A2(n132), .ZN(n4071) );
  OR2_X1 U625 ( .A1(n3984), .A2(n3983), .ZN(n4072) );
  NAND2_X2 U626 ( .A1(n4175), .A2(n1631), .ZN(n4177) );
  INV_X2 U627 ( .A(n4073), .ZN(n1636) );
  NAND2_X2 U631 ( .A1(n4003), .A2(n3978), .ZN(n4073) );
  NAND2_X2 U632 ( .A1(n1789), .A2(n1632), .ZN(n2118) );
  OAI21_X2 U639 ( .B1(n720), .B2(n719), .A(n718), .ZN(n1789) );
  INV_X1 U641 ( .A(n999), .ZN(n4074) );
  NAND2_X2 U644 ( .A1(n1478), .A2(n1336), .ZN(n4075) );
  NAND2_X2 U656 ( .A1(n1478), .A2(n1336), .ZN(n3460) );
  AND2_X2 U657 ( .A1(b[2]), .A2(n2506), .ZN(n1336) );
  NAND2_X4 U672 ( .A1(n4102), .A2(n307), .ZN(n1232) );
  NAND2_X1 U675 ( .A1(n3177), .A2(n3534), .ZN(n2870) );
  NAND2_X4 U687 ( .A1(n3607), .A2(n3608), .ZN(n3978) );
  INV_X4 U690 ( .A(n1795), .ZN(n681) );
  NAND2_X2 U691 ( .A1(n4084), .A2(n4081), .ZN(n4076) );
  INV_X1 U696 ( .A(n2961), .ZN(n2276) );
  NOR2_X2 U700 ( .A1(n1015), .A2(n2957), .ZN(n2961) );
  INV_X1 U703 ( .A(n2288), .ZN(n3105) );
  NAND2_X1 U704 ( .A1(n3063), .A2(n3064), .ZN(n3084) );
  NAND2_X2 U706 ( .A1(n4104), .A2(n4103), .ZN(n4077) );
  NAND2_X1 U708 ( .A1(a[23]), .A2(n1913), .ZN(n1228) );
  INV_X4 U709 ( .A(n3097), .ZN(n1577) );
  INV_X2 U719 ( .A(n1540), .ZN(n4078) );
  INV_X2 U720 ( .A(n4078), .ZN(n4079) );
  INV_X1 U721 ( .A(n3050), .ZN(n1531) );
  NAND3_X2 U725 ( .A1(n4139), .A2(n400), .A3(n2852), .ZN(n2197) );
  INV_X4 U727 ( .A(n1165), .ZN(n976) );
  NAND2_X2 U729 ( .A1(n666), .A2(n1965), .ZN(n161) );
  NAND2_X2 U730 ( .A1(n1970), .A2(n1805), .ZN(n666) );
  NAND2_X2 U733 ( .A1(n2950), .A2(n2949), .ZN(n1810) );
  NAND2_X2 U738 ( .A1(n976), .A2(n2933), .ZN(n2950) );
  NAND2_X2 U739 ( .A1(n2275), .A2(n2963), .ZN(n198) );
  NAND2_X2 U742 ( .A1(n2140), .A2(n2141), .ZN(n2275) );
  NAND2_X2 U763 ( .A1(n3272), .A2(n69), .ZN(n322) );
  NAND2_X2 U767 ( .A1(n324), .A2(n2564), .ZN(n3272) );
  NAND3_X2 U777 ( .A1(n1139), .A2(n2197), .A3(n2116), .ZN(n2114) );
  NAND2_X2 U778 ( .A1(n2054), .A2(n2055), .ZN(n3104) );
  OAI21_X2 U782 ( .B1(n103), .B2(n2377), .A(n2226), .ZN(n2054) );
  AOI22_X2 U783 ( .A1(n521), .A2(n4080), .B1(n520), .B2(n3969), .ZN(n3734) );
  AOI22_X2 U788 ( .A1(n2344), .A2(n2343), .B1(n2342), .B2(n59), .ZN(n4080) );
  NAND2_X2 U790 ( .A1(n2188), .A2(n3092), .ZN(n3097) );
  NAND2_X2 U791 ( .A1(n1217), .A2(n3208), .ZN(n2241) );
  INV_X2 U805 ( .A(n775), .ZN(n774) );
  NAND2_X2 U815 ( .A1(n776), .A2(n777), .ZN(n775) );
  OAI21_X2 U826 ( .B1(n2851), .B2(n2850), .A(n2853), .ZN(n400) );
  NAND3_X2 U828 ( .A1(n2287), .A2(n2175), .A3(n2176), .ZN(n1960) );
  NAND2_X2 U832 ( .A1(n4084), .A2(n4081), .ZN(n3234) );
  NAND2_X2 U839 ( .A1(n4083), .A2(n4082), .ZN(n4081) );
  INV_X2 U851 ( .A(n2029), .ZN(n4083) );
  NAND2_X2 U871 ( .A1(n3231), .A2(n3230), .ZN(n4084) );
  NAND2_X2 U884 ( .A1(n2048), .A2(n2218), .ZN(n957) );
  NAND3_X1 U887 ( .A1(n2220), .A2(n2219), .A3(n2789), .ZN(n2218) );
  NAND2_X2 U916 ( .A1(n3431), .A2(n1554), .ZN(n2287) );
  NOR2_X2 U917 ( .A1(n1123), .A2(n2114), .ZN(n1866) );
  INV_X4 U920 ( .A(n1917), .ZN(n1123) );
  NAND2_X2 U921 ( .A1(n4104), .A2(n4103), .ZN(n1917) );
  NAND2_X2 U926 ( .A1(n1810), .A2(n1809), .ZN(n1565) );
  NAND2_X1 U931 ( .A1(n3206), .A2(a[23]), .ZN(n2458) );
  NAND2_X4 U937 ( .A1(n2199), .A2(n3027), .ZN(n3206) );
  NAND3_X2 U938 ( .A1(n2140), .A2(n2963), .A3(n2141), .ZN(n1959) );
  NAND2_X2 U939 ( .A1(n2015), .A2(n2954), .ZN(n2140) );
  BUF_X4 U945 ( .A(n85), .Z(n4085) );
  INV_X4 U952 ( .A(n4086), .ZN(n2013) );
  NOR2_X2 U964 ( .A1(n532), .A2(n531), .ZN(n4086) );
  NAND2_X2 U965 ( .A1(n3915), .A2(n3715), .ZN(n3729) );
  NAND2_X4 U967 ( .A1(n951), .A2(n2679), .ZN(n3915) );
  INV_X2 U971 ( .A(n4087), .ZN(n4198) );
  NAND2_X2 U977 ( .A1(n2931), .A2(n2930), .ZN(n4087) );
  NAND2_X2 U978 ( .A1(n2078), .A2(n4088), .ZN(n950) );
  OAI22_X2 U999 ( .A1(n3644), .A2(n2271), .B1(n4090), .B2(n1705), .ZN(n245) );
  XNOR2_X2 U1003 ( .A(n3389), .B(n3010), .ZN(n4090) );
  NAND2_X2 U1006 ( .A1(n1994), .A2(n1992), .ZN(n1723) );
  NAND2_X2 U1010 ( .A1(n1724), .A2(n1725), .ZN(n1994) );
  NAND2_X2 U1013 ( .A1(n793), .A2(n400), .ZN(n792) );
  NOR2_X2 U1014 ( .A1(n1961), .A2(n2043), .ZN(n2970) );
  NAND2_X2 U1017 ( .A1(n1372), .A2(n1373), .ZN(n1133) );
  NAND2_X2 U1023 ( .A1(n2603), .A2(n2605), .ZN(n1372) );
  XNOR2_X2 U1035 ( .A(n4091), .B(n2480), .ZN(n932) );
  NAND2_X2 U1046 ( .A1(n1431), .A2(n1430), .ZN(n4091) );
  NAND2_X2 U1048 ( .A1(n433), .A2(n2772), .ZN(n1587) );
  NAND2_X2 U1054 ( .A1(n838), .A2(n837), .ZN(n433) );
  NAND2_X2 U1073 ( .A1(n4092), .A2(n3079), .ZN(n177) );
  INV_X2 U1080 ( .A(n3302), .ZN(n4092) );
  NAND2_X2 U1082 ( .A1(n3301), .A2(n3300), .ZN(n3302) );
  NOR2_X1 U1090 ( .A1(n3535), .A2(n3505), .ZN(n3528) );
  NAND2_X2 U1093 ( .A1(n3526), .A2(n1670), .ZN(n1669) );
  NOR2_X2 U1104 ( .A1(n1142), .A2(n1145), .ZN(n3526) );
  INV_X2 U1107 ( .A(n1180), .ZN(n4093) );
  NAND2_X2 U1110 ( .A1(n2513), .A2(n4093), .ZN(n128) );
  NAND2_X2 U1112 ( .A1(n4094), .A2(n1344), .ZN(n2186) );
  NAND2_X2 U1120 ( .A1(n1343), .A2(n3190), .ZN(n4094) );
  NOR2_X2 U1121 ( .A1(b[2]), .A2(n2506), .ZN(n4154) );
  NAND2_X2 U1122 ( .A1(n4095), .A2(n2857), .ZN(n1553) );
  NAND2_X2 U1123 ( .A1(n243), .A2(n245), .ZN(n2857) );
  NAND2_X2 U1132 ( .A1(n9), .A2(n4131), .ZN(n4095) );
  NOR2_X1 U1141 ( .A1(n2395), .A2(n1022), .ZN(n2297) );
  NAND3_X2 U1142 ( .A1(n398), .A2(n4180), .A3(n1856), .ZN(n2395) );
  NAND2_X2 U1152 ( .A1(n3873), .A2(n3915), .ZN(n3878) );
  INV_X8 U1164 ( .A(n3915), .ZN(n3924) );
  INV_X4 U1168 ( .A(n3535), .ZN(n3495) );
  NAND2_X2 U1169 ( .A1(n4096), .A2(n3246), .ZN(n1073) );
  INV_X2 U1172 ( .A(n1647), .ZN(n4096) );
  NAND2_X2 U1183 ( .A1(n1521), .A2(n1520), .ZN(n1647) );
  NOR2_X2 U1187 ( .A1(n4156), .A2(n1907), .ZN(n2010) );
  NOR2_X2 U1192 ( .A1(n2103), .A2(n2104), .ZN(n4156) );
  NAND2_X2 U1193 ( .A1(n3119), .A2(n2941), .ZN(n4126) );
  NOR2_X2 U1194 ( .A1(n763), .A2(n1604), .ZN(n1603) );
  NAND2_X2 U1196 ( .A1(n730), .A2(n729), .ZN(n763) );
  OR2_X2 U1201 ( .A1(n3310), .A2(a[9]), .ZN(n1978) );
  NAND2_X2 U1203 ( .A1(n4125), .A2(n4124), .ZN(n1907) );
  INV_X4 U1211 ( .A(n1202), .ZN(n4008) );
  NAND2_X2 U1212 ( .A1(n3736), .A2(n3737), .ZN(n1202) );
  AOI22_X2 U1219 ( .A1(n4097), .A2(n3999), .B1(n931), .B2(n3937), .ZN(n3942)
         );
  NOR2_X4 U1221 ( .A1(n4018), .A2(n3936), .ZN(n4097) );
  OAI21_X2 U1228 ( .B1(n2350), .B2(n2353), .A(n24), .ZN(n3300) );
  OR2_X2 U1235 ( .A1(n2998), .A2(n1600), .ZN(n3075) );
  NAND3_X2 U1257 ( .A1(n2093), .A2(n2352), .A3(n2351), .ZN(n3301) );
  NOR2_X4 U1259 ( .A1(n4098), .A2(n3448), .ZN(n3557) );
  NOR2_X2 U1261 ( .A1(n1650), .A2(n3446), .ZN(n4098) );
  NOR2_X2 U1262 ( .A1(n2165), .A2(n2924), .ZN(n4099) );
  INV_X1 U1263 ( .A(n3866), .ZN(n3659) );
  NAND2_X2 U1267 ( .A1(n3579), .A2(n3580), .ZN(n3866) );
  NAND2_X2 U1268 ( .A1(n1734), .A2(n1733), .ZN(n1379) );
  OAI21_X2 U1269 ( .B1(n1198), .B2(n1685), .A(n2905), .ZN(n1734) );
  INV_X2 U1270 ( .A(n2815), .ZN(n1537) );
  NAND2_X2 U1275 ( .A1(n231), .A2(n1163), .ZN(n2815) );
  INV_X4 U1279 ( .A(n2937), .ZN(n103) );
  NAND2_X2 U1282 ( .A1(n1504), .A2(n1503), .ZN(n1165) );
  NAND2_X2 U1283 ( .A1(n717), .A2(n716), .ZN(n1632) );
  NAND3_X2 U1291 ( .A1(n1076), .A2(n1959), .A3(n2965), .ZN(n1503) );
  INV_X2 U1292 ( .A(n1169), .ZN(n1354) );
  NAND2_X2 U1293 ( .A1(n4205), .A2(n322), .ZN(n1169) );
  NAND2_X2 U1294 ( .A1(n844), .A2(n845), .ZN(n2625) );
  NAND2_X2 U1301 ( .A1(n4100), .A2(n1012), .ZN(n1010) );
  NOR2_X2 U1305 ( .A1(n2277), .A2(n927), .ZN(n4100) );
  NAND3_X2 U1307 ( .A1(n2231), .A2(n2234), .A3(n2233), .ZN(n1795) );
  NAND2_X2 U1308 ( .A1(n1881), .A2(n2029), .ZN(n752) );
  INV_X1 U1310 ( .A(n3505), .ZN(n4101) );
  NOR2_X1 U1311 ( .A1(n3532), .A2(n4101), .ZN(n455) );
  NAND2_X2 U1315 ( .A1(n1390), .A2(n1389), .ZN(n4102) );
  NOR2_X2 U1316 ( .A1(n4024), .A2(n3612), .ZN(n3714) );
  NAND2_X2 U1317 ( .A1(n3611), .A2(n1848), .ZN(n4024) );
  NAND3_X2 U1326 ( .A1(n2894), .A2(n1915), .A3(n1916), .ZN(n4103) );
  OAI21_X2 U1338 ( .B1(n1122), .B2(n1280), .A(n1914), .ZN(n4104) );
  NAND2_X2 U1366 ( .A1(n1936), .A2(n4105), .ZN(n1022) );
  NAND3_X1 U1372 ( .A1(n1474), .A2(n3021), .A3(n3022), .ZN(n4105) );
  NAND2_X2 U1374 ( .A1(n834), .A2(n4106), .ZN(n2979) );
  NAND2_X2 U1379 ( .A1(n4129), .A2(n3139), .ZN(n4106) );
  INV_X4 U1392 ( .A(n2925), .ZN(n1610) );
  NAND2_X2 U1401 ( .A1(n2198), .A2(n2407), .ZN(n1358) );
  INV_X4 U1402 ( .A(n4107), .ZN(n1575) );
  NOR2_X4 U1411 ( .A1(n2285), .A2(n2994), .ZN(n4107) );
  NAND2_X2 U1414 ( .A1(n4108), .A2(n1109), .ZN(n430) );
  NAND2_X2 U1418 ( .A1(n1417), .A2(n1416), .ZN(n4108) );
  NAND2_X2 U1437 ( .A1(n116), .A2(n2846), .ZN(n2937) );
  NAND2_X2 U1462 ( .A1(n4110), .A2(n4109), .ZN(n1910) );
  INV_X2 U1465 ( .A(n2104), .ZN(n4109) );
  INV_X2 U1508 ( .A(n2103), .ZN(n4110) );
  NAND2_X2 U1517 ( .A1(n2384), .A2(n37), .ZN(n1699) );
  NOR2_X2 U1518 ( .A1(n4112), .A2(n4111), .ZN(n547) );
  NAND2_X2 U1523 ( .A1(n1624), .A2(n1625), .ZN(n4111) );
  INV_X2 U1527 ( .A(n1957), .ZN(n4112) );
  NAND2_X2 U1528 ( .A1(n4114), .A2(n4113), .ZN(n1594) );
  INV_X2 U1533 ( .A(n675), .ZN(n4113) );
  INV_X2 U1545 ( .A(n2147), .ZN(n4114) );
  XNOR2_X2 U1574 ( .A(n4117), .B(n3385), .ZN(n3387) );
  NAND3_X2 U1575 ( .A1(n301), .A2(n300), .A3(n3384), .ZN(n4117) );
  NAND2_X2 U1613 ( .A1(n1160), .A2(n817), .ZN(n1605) );
  NAND2_X2 U1631 ( .A1(n118), .A2(n119), .ZN(n1160) );
  NAND2_X2 U1635 ( .A1(n3239), .A2(n3238), .ZN(n3277) );
  INV_X4 U1639 ( .A(n4118), .ZN(n387) );
  NOR2_X2 U1659 ( .A1(n3255), .A2(n540), .ZN(n4118) );
  NAND2_X2 U1673 ( .A1(n1902), .A2(n1899), .ZN(n3607) );
  NAND3_X2 U1733 ( .A1(n1901), .A2(n3267), .A3(n1900), .ZN(n1899) );
  OAI21_X2 U1734 ( .B1(n1903), .B2(n2331), .A(n3268), .ZN(n1902) );
  NAND3_X2 U1751 ( .A1(n3638), .A2(n3637), .A3(n3864), .ZN(n855) );
  NAND2_X4 U1766 ( .A1(n337), .A2(n4119), .ZN(n3573) );
  NAND3_X2 U1776 ( .A1(n336), .A2(n3381), .A3(n1878), .ZN(n4119) );
  NOR3_X2 U1808 ( .A1(n2765), .A2(n2767), .A3(n4120), .ZN(n1790) );
  NOR3_X2 U1817 ( .A1(n4208), .A2(n2764), .A3(n2760), .ZN(n4120) );
  NAND2_X2 U1820 ( .A1(n1335), .A2(n1334), .ZN(n2564) );
  NAND2_X2 U1831 ( .A1(n3066), .A2(n2556), .ZN(n2193) );
  NOR2_X2 U1845 ( .A1(n2561), .A2(n2560), .ZN(n3269) );
  AOI21_X2 U1849 ( .B1(n370), .B2(n3292), .A(n369), .ZN(n2560) );
  OAI22_X2 U1859 ( .A1(n1227), .A2(a[25]), .B1(n1478), .B2(n2434), .ZN(n1687)
         );
  NAND2_X2 U1860 ( .A1(n4121), .A2(n1296), .ZN(n2774) );
  NAND2_X2 U1861 ( .A1(n1294), .A2(n1295), .ZN(n4121) );
  INV_X4 U1887 ( .A(n4122), .ZN(n3249) );
  NOR2_X2 U1889 ( .A1(n3294), .A2(n811), .ZN(n4122) );
  NAND2_X2 U1902 ( .A1(n1587), .A2(n4123), .ZN(n2064) );
  NAND3_X1 U1903 ( .A1(n348), .A2(n837), .A3(n838), .ZN(n4123) );
  NAND2_X1 U1937 ( .A1(n4035), .A2(n1360), .ZN(n50) );
  INV_X2 U1938 ( .A(n607), .ZN(n4124) );
  NAND2_X2 U1944 ( .A1(n608), .A2(n3199), .ZN(n4125) );
  NAND2_X2 U1957 ( .A1(n2352), .A2(n2351), .ZN(n2350) );
  NAND2_X2 U1958 ( .A1(n86), .A2(n2356), .ZN(n2352) );
  NAND2_X2 U1982 ( .A1(n435), .A2(n2306), .ZN(n3732) );
  INV_X2 U2024 ( .A(n3371), .ZN(n1214) );
  XNOR2_X2 U2039 ( .A(n691), .B(n690), .ZN(n3371) );
  INV_X2 U2044 ( .A(n2167), .ZN(n1436) );
  NAND2_X2 U2051 ( .A1(n507), .A2(n506), .ZN(n2167) );
  NAND2_X2 U2054 ( .A1(n4126), .A2(n1327), .ZN(n2451) );
  NOR2_X2 U2066 ( .A1(n2509), .A2(n2508), .ZN(n2511) );
  NOR2_X2 U2079 ( .A1(n2417), .A2(n2418), .ZN(n2509) );
  NAND3_X2 U2080 ( .A1(n4128), .A2(n1228), .A3(n57), .ZN(n4127) );
  NAND2_X2 U2100 ( .A1(n1227), .A2(n45), .ZN(n4128) );
  INV_X1 U2113 ( .A(n1449), .ZN(n4129) );
  NAND2_X2 U2125 ( .A1(n4130), .A2(n4209), .ZN(n3366) );
  NOR2_X2 U2127 ( .A1(n1029), .A2(n3041), .ZN(n4130) );
  INV_X2 U2134 ( .A(n245), .ZN(n4131) );
  NAND2_X2 U2139 ( .A1(n1371), .A2(n3700), .ZN(n3702) );
  NAND2_X2 U2140 ( .A1(n2247), .A2(n3990), .ZN(n1371) );
  INV_X2 U2150 ( .A(n2538), .ZN(n3210) );
  XNOR2_X1 U2151 ( .A(n1323), .B(a[15]), .ZN(n2538) );
  NAND2_X2 U2156 ( .A1(n1840), .A2(n4132), .ZN(n2375) );
  NOR2_X2 U2158 ( .A1(n2948), .A2(n2946), .ZN(n4132) );
  OAI21_X2 U2173 ( .B1(n4013), .B2(n4015), .A(n4133), .ZN(n4014) );
  AOI22_X2 U2176 ( .A1(n237), .A2(n678), .B1(n4012), .B2(n679), .ZN(n4133) );
  NAND2_X2 U2180 ( .A1(n1659), .A2(a[20]), .ZN(n3110) );
  NAND2_X2 U2199 ( .A1(n2657), .A2(n2658), .ZN(n2758) );
  NAND2_X2 U2201 ( .A1(n2867), .A2(n2866), .ZN(n1480) );
  NAND3_X2 U2207 ( .A1(n769), .A2(n4134), .A3(n1283), .ZN(n766) );
  INV_X2 U2208 ( .A(n885), .ZN(n4134) );
  NOR2_X2 U2214 ( .A1(n3292), .A2(n3291), .ZN(n885) );
  NAND2_X2 U2215 ( .A1(n4135), .A2(n1592), .ZN(n887) );
  INV_X2 U2216 ( .A(n2547), .ZN(n4135) );
  NAND2_X2 U2222 ( .A1(n2523), .A2(n2522), .ZN(n2547) );
  NAND2_X2 U2223 ( .A1(n2383), .A2(n2087), .ZN(n110) );
  NOR2_X4 U2226 ( .A1(n4136), .A2(n3002), .ZN(n3053) );
  NAND2_X2 U2229 ( .A1(n1731), .A2(n1732), .ZN(n4136) );
  NAND2_X2 U2233 ( .A1(n111), .A2(n93), .ZN(n1918) );
  NAND2_X2 U2234 ( .A1(n2139), .A2(n2925), .ZN(n2963) );
  INV_X2 U2236 ( .A(n4137), .ZN(n1086) );
  NOR2_X2 U2239 ( .A1(n3239), .A2(n3238), .ZN(n4137) );
  NAND2_X2 U2244 ( .A1(n4138), .A2(n1760), .ZN(n312) );
  NAND3_X2 U2252 ( .A1(n1932), .A2(n402), .A3(n2888), .ZN(n4138) );
  INV_X4 U2263 ( .A(n3026), .ZN(n4155) );
  AOI21_X1 U2265 ( .B1(n3217), .B2(n1863), .A(n1738), .ZN(n1176) );
  NAND2_X2 U2266 ( .A1(n672), .A2(n671), .ZN(n1683) );
  INV_X2 U2277 ( .A(n4027), .ZN(n1571) );
  INV_X1 U2282 ( .A(n536), .ZN(n535) );
  OAI21_X1 U2293 ( .B1(n536), .B2(n284), .A(n3960), .ZN(n533) );
  AOI21_X2 U2302 ( .B1(n3444), .B2(n924), .A(n3443), .ZN(n2180) );
  NAND2_X2 U2308 ( .A1(n256), .A2(n255), .ZN(n4139) );
  NAND2_X2 U2309 ( .A1(n1585), .A2(n3350), .ZN(n4140) );
  NAND2_X2 U2310 ( .A1(n1585), .A2(n3350), .ZN(n822) );
  NOR2_X2 U2312 ( .A1(n749), .A2(n750), .ZN(n2477) );
  NAND2_X1 U2323 ( .A1(n2477), .A2(n737), .ZN(n1406) );
  INV_X1 U2330 ( .A(n2477), .ZN(n1140) );
  NAND2_X2 U2332 ( .A1(n736), .A2(n2477), .ZN(n733) );
  AOI21_X1 U2335 ( .B1(n1649), .B2(n3407), .A(n2322), .ZN(n1025) );
  NAND2_X1 U2336 ( .A1(n2318), .A2(n2940), .ZN(n1046) );
  NAND2_X2 U2341 ( .A1(n1416), .A2(n1417), .ZN(n1110) );
  INV_X2 U2349 ( .A(n1605), .ZN(n3318) );
  NAND2_X1 U2361 ( .A1(n3980), .A2(n3979), .ZN(n1524) );
  NAND2_X1 U2362 ( .A1(n3977), .A2(n3759), .ZN(n3758) );
  INV_X1 U2365 ( .A(n3977), .ZN(n4189) );
  NAND2_X2 U2371 ( .A1(n133), .A2(n132), .ZN(n4141) );
  NAND2_X2 U2376 ( .A1(n109), .A2(n4071), .ZN(n4142) );
  INV_X2 U2384 ( .A(n1141), .ZN(n1258) );
  AOI22_X2 U2386 ( .A1(n3435), .A2(n3395), .B1(n2182), .B2(n3394), .ZN(n4143)
         );
  NAND2_X1 U2387 ( .A1(n598), .A2(n3397), .ZN(n4146) );
  NAND2_X2 U2408 ( .A1(n4146), .A2(n4147), .ZN(n3444) );
  NOR2_X1 U2426 ( .A1(n3439), .A2(n3444), .ZN(n221) );
  NOR2_X1 U2436 ( .A1(n3444), .A2(n924), .ZN(n2179) );
  INV_X1 U2437 ( .A(n3444), .ZN(n590) );
  OAI21_X1 U2438 ( .B1(n2935), .B2(n2948), .A(n2946), .ZN(n2373) );
  OAI21_X1 U2440 ( .B1(n2935), .B2(n2948), .A(n2946), .ZN(n2370) );
  INV_X2 U2454 ( .A(n3702), .ZN(n2062) );
  INV_X1 U2461 ( .A(n2248), .ZN(n3988) );
  AND2_X2 U2463 ( .A1(n2740), .A2(n2741), .ZN(n3076) );
  INV_X2 U2464 ( .A(n2985), .ZN(n1455) );
  INV_X2 U2495 ( .A(n249), .ZN(n4149) );
  NAND2_X1 U2497 ( .A1(n550), .A2(n549), .ZN(n4150) );
  INV_X2 U2500 ( .A(n3541), .ZN(n74) );
  AOI21_X1 U2505 ( .B1(n1618), .B2(n4010), .A(n4009), .ZN(n678) );
  NOR2_X4 U2516 ( .A1(n382), .A2(n381), .ZN(n719) );
  AOI22_X1 U2517 ( .A1(n2027), .A2(n2356), .B1(n4044), .B2(n3034), .ZN(n1860)
         );
  NAND2_X1 U2522 ( .A1(n3034), .A2(n94), .ZN(n1981) );
  NOR2_X1 U2524 ( .A1(n3176), .A2(n3109), .ZN(n1340) );
  NAND2_X2 U2528 ( .A1(n1639), .A2(n1447), .ZN(n2237) );
  NAND2_X2 U2538 ( .A1(n705), .A2(n64), .ZN(n4151) );
  AND3_X1 U2539 ( .A1(n2281), .A2(n1701), .A3(n1232), .ZN(n4152) );
  INV_X8 U2540 ( .A(n1510), .ZN(n1639) );
  INV_X1 U2547 ( .A(n2423), .ZN(n2301) );
  NAND2_X4 U2560 ( .A1(n2209), .A2(n2125), .ZN(n194) );
  NOR2_X2 U2564 ( .A1(n2112), .A2(n19), .ZN(n1141) );
  INV_X1 U2581 ( .A(n2112), .ZN(n265) );
  NAND2_X1 U2598 ( .A1(n19), .A2(n2112), .ZN(n1259) );
  NAND3_X2 U2607 ( .A1(n3516), .A2(n3515), .A3(n3535), .ZN(n3519) );
  NOR2_X1 U2610 ( .A1(n3168), .A2(n3169), .ZN(n4153) );
  NOR2_X2 U2617 ( .A1(n3168), .A2(n3169), .ZN(n1786) );
  NAND2_X2 U2618 ( .A1(n2282), .A2(n1281), .ZN(n1474) );
  NAND2_X2 U2620 ( .A1(n4154), .A2(n2556), .ZN(n1928) );
  INV_X4 U2621 ( .A(n257), .ZN(n256) );
  XOR2_X1 U2624 ( .A(n4023), .B(n4157), .Z(\d[22]_BAR ) );
  OR2_X1 U2637 ( .A1(n3961), .A2(n1787), .ZN(n4157) );
  INV_X8 U2640 ( .A(n2506), .ZN(n3065) );
  INV_X1 U2641 ( .A(n1940), .ZN(n1005) );
  INV_X1 U2643 ( .A(n2043), .ZN(n1053) );
  NAND2_X1 U2644 ( .A1(n289), .A2(n285), .ZN(n4158) );
  INV_X1 U2655 ( .A(n1414), .ZN(n4159) );
  INV_X1 U2658 ( .A(n3398), .ZN(n1414) );
  NAND2_X1 U2663 ( .A1(n1862), .A2(n3407), .ZN(n421) );
  NAND2_X1 U2675 ( .A1(n1862), .A2(n90), .ZN(n180) );
  NAND2_X1 U2676 ( .A1(n1862), .A2(n37), .ZN(n2176) );
  NAND2_X1 U2681 ( .A1(n1694), .A2(n1693), .ZN(n3404) );
  NOR2_X1 U2689 ( .A1(n82), .A2(n3535), .ZN(n779) );
  AND2_X1 U2690 ( .A1(n4038), .A2(n421), .ZN(n49) );
  NAND2_X1 U2691 ( .A1(n180), .A2(n179), .ZN(n178) );
  NAND3_X1 U2694 ( .A1(n3089), .A2(n3088), .A3(n431), .ZN(n3091) );
  NOR2_X1 U2696 ( .A1(n634), .A2(n633), .ZN(n4161) );
  INV_X2 U2700 ( .A(n2647), .ZN(n2651) );
  INV_X4 U2715 ( .A(n1997), .ZN(n1138) );
  NAND2_X1 U2716 ( .A1(n619), .A2(n2961), .ZN(n4164) );
  NAND2_X2 U2721 ( .A1(n4164), .A2(n4165), .ZN(n1569) );
  NAND2_X2 U2729 ( .A1(n2139), .A2(n1610), .ZN(n4166) );
  NAND2_X2 U2730 ( .A1(n2139), .A2(n1610), .ZN(n1612) );
  NAND2_X1 U2732 ( .A1(n4075), .A2(a[23]), .ZN(n280) );
  XNOR2_X1 U2736 ( .A(n3537), .B(n4167), .ZN(n3539) );
  INV_X1 U2756 ( .A(n3552), .ZN(n4167) );
  INV_X1 U2765 ( .A(n3537), .ZN(n3547) );
  NAND2_X2 U2780 ( .A1(n2540), .A2(n2539), .ZN(n3251) );
  NAND2_X1 U2783 ( .A1(n599), .A2(n1578), .ZN(n3745) );
  INV_X4 U2789 ( .A(n2555), .ZN(n2122) );
  NAND2_X1 U2793 ( .A1(n3086), .A2(n65), .ZN(n170) );
  INV_X1 U2795 ( .A(n3435), .ZN(n1548) );
  AND2_X2 U2800 ( .A1(n1532), .A2(n1533), .ZN(n446) );
  NAND2_X1 U2820 ( .A1(n1532), .A2(n1533), .ZN(n1324) );
  INV_X2 U2827 ( .A(n2382), .ZN(n2441) );
  INV_X4 U2845 ( .A(n3940), .ZN(n3999) );
  OAI21_X2 U2859 ( .B1(n459), .B2(n1762), .A(n3010), .ZN(n1861) );
  NAND2_X1 U2862 ( .A1(n1626), .A2(n1630), .ZN(n3280) );
  NAND2_X1 U2868 ( .A1(n2041), .A2(n2042), .ZN(n610) );
  NOR2_X4 U2870 ( .A1(n3305), .A2(n3304), .ZN(n3333) );
  INV_X2 U2876 ( .A(n2976), .ZN(n4168) );
  INV_X2 U2877 ( .A(n4168), .ZN(n4169) );
  NAND2_X1 U2901 ( .A1(n3710), .A2(n1586), .ZN(n3628) );
  NAND2_X1 U2902 ( .A1(n820), .A2(n3710), .ZN(n2290) );
  NAND2_X1 U2910 ( .A1(n3685), .A2(n3710), .ZN(n3677) );
  INV_X4 U2915 ( .A(n1101), .ZN(n1585) );
  NAND2_X4 U2918 ( .A1(n387), .A2(n386), .ZN(n3257) );
  OAI21_X2 U2923 ( .B1(n2007), .B2(n3564), .A(n3567), .ZN(n1395) );
  NAND2_X2 U2952 ( .A1(n1441), .A2(n2559), .ZN(n1442) );
  NOR2_X2 U2959 ( .A1(n856), .A2(n3619), .ZN(n3638) );
  INV_X2 U2972 ( .A(n2772), .ZN(n348) );
  MUX2_X1 U2988 ( .A(n1303), .B(n3204), .S(a[20]), .Z(n2640) );
  MUX2_X1 U2989 ( .A(n1303), .B(n3204), .S(a[17]), .Z(n2466) );
  OR2_X2 U2992 ( .A1(n1303), .A2(a[3]), .ZN(n17) );
  NOR2_X2 U2993 ( .A1(n1303), .A2(n93), .ZN(n615) );
  INV_X2 U3003 ( .A(n3352), .ZN(n1240) );
  NAND2_X1 U3005 ( .A1(n3353), .A2(n3352), .ZN(n1241) );
  NAND2_X2 U3008 ( .A1(b[3]), .A2(n4171), .ZN(n4172) );
  NAND2_X2 U3009 ( .A1(n4170), .A2(b[4]), .ZN(n4173) );
  NAND2_X2 U3014 ( .A1(n4172), .A2(n4173), .ZN(n2382) );
  INV_X2 U3016 ( .A(b[3]), .ZN(n4170) );
  INV_X2 U3018 ( .A(b[4]), .ZN(n4171) );
  OAI21_X1 U3023 ( .B1(n84), .B2(n1784), .A(n2156), .ZN(n498) );
  NOR2_X4 U3031 ( .A1(n1600), .A2(b[11]), .ZN(n2742) );
  NOR2_X1 U3041 ( .A1(n2401), .A2(n432), .ZN(n2313) );
  NAND2_X2 U3050 ( .A1(n1882), .A2(n650), .ZN(n4174) );
  NOR2_X4 U3070 ( .A1(n1745), .A2(n3947), .ZN(n3572) );
  NAND2_X2 U3078 ( .A1(n2186), .A2(n3192), .ZN(n11) );
  NAND3_X1 U3081 ( .A1(n1208), .A2(n1630), .A3(n3277), .ZN(n4202) );
  NAND2_X2 U3130 ( .A1(n707), .A2(n709), .ZN(n706) );
  NAND2_X4 U3133 ( .A1(n1765), .A2(n1317), .ZN(n3305) );
  INV_X2 U3140 ( .A(n3966), .ZN(n3967) );
  NAND2_X1 U3141 ( .A1(n3087), .A2(n2992), .ZN(n303) );
  NAND2_X1 U3151 ( .A1(n3286), .A2(n3271), .ZN(n4176) );
  NAND2_X2 U3152 ( .A1(n4176), .A2(n4177), .ZN(n1988) );
  INV_X2 U3158 ( .A(n3286), .ZN(n4175) );
  NAND2_X2 U3167 ( .A1(n2919), .A2(n775), .ZN(n405) );
  INV_X2 U3169 ( .A(n842), .ZN(n2656) );
  NOR2_X4 U3170 ( .A1(n3573), .A2(n3574), .ZN(n3612) );
  INV_X2 U3173 ( .A(n1916), .ZN(n1122) );
  NOR2_X4 U3174 ( .A1(n151), .A2(n2214), .ZN(n1914) );
  NOR2_X1 U3175 ( .A1(n3702), .A2(n3701), .ZN(n3704) );
  NAND2_X1 U3178 ( .A1(n544), .A2(n2512), .ZN(n543) );
  AOI21_X2 U3180 ( .B1(n3028), .B2(n3029), .A(n3030), .ZN(n4178) );
  INV_X2 U3181 ( .A(n3089), .ZN(n4179) );
  INV_X1 U3184 ( .A(n3290), .ZN(n424) );
  NAND2_X2 U3214 ( .A1(n773), .A2(n774), .ZN(n406) );
  NOR2_X4 U3224 ( .A1(b[7]), .A2(b[8]), .ZN(n2689) );
  INV_X4 U3227 ( .A(n3269), .ZN(n377) );
  NAND2_X1 U3234 ( .A1(n1737), .A2(n3988), .ZN(n3940) );
  NAND2_X1 U3244 ( .A1(n3089), .A2(n1124), .ZN(n4180) );
  NAND2_X2 U3245 ( .A1(n2135), .A2(n2134), .ZN(n4181) );
  NAND2_X1 U3248 ( .A1(n3057), .A2(n1313), .ZN(n3055) );
  NOR2_X1 U3252 ( .A1(n3915), .A2(n3628), .ZN(n3631) );
  NOR2_X1 U3257 ( .A1(n3915), .A2(n3677), .ZN(n3695) );
  NAND2_X2 U3259 ( .A1(n3266), .A2(n2294), .ZN(n3737) );
  INV_X4 U3265 ( .A(n194), .ZN(n2068) );
  NAND2_X2 U3266 ( .A1(n3180), .A2(n3185), .ZN(n1282) );
  INV_X2 U3283 ( .A(n3192), .ZN(n1466) );
  NAND2_X4 U3285 ( .A1(n1300), .A2(n2947), .ZN(n1840) );
  NAND2_X4 U3301 ( .A1(n404), .A2(n403), .ZN(n2947) );
  INV_X2 U3306 ( .A(n1685), .ZN(n2293) );
  NOR2_X1 U3313 ( .A1(n4181), .A2(n142), .ZN(n4182) );
  AOI22_X2 U3325 ( .A1(n3034), .A2(n3413), .B1(n3407), .B2(n3177), .ZN(n2143)
         );
  NAND2_X1 U3328 ( .A1(n169), .A2(n3092), .ZN(n506) );
  NAND3_X1 U3331 ( .A1(n3070), .A2(n1890), .A3(n2193), .ZN(n1370) );
  NAND2_X1 U3351 ( .A1(n2174), .A2(b[2]), .ZN(n4184) );
  NAND2_X2 U3358 ( .A1(n4183), .A2(n3066), .ZN(n4185) );
  NAND2_X4 U3362 ( .A1(n4184), .A2(n4185), .ZN(n1898) );
  INV_X2 U3363 ( .A(n2174), .ZN(n4183) );
  NOR3_X2 U3370 ( .A1(n3747), .A2(n1497), .A3(n2011), .ZN(n522) );
  NAND3_X2 U3372 ( .A1(n1908), .A2(n1909), .A3(n1906), .ZN(n2209) );
  NAND2_X2 U3374 ( .A1(n3758), .A2(n4187), .ZN(\d[19] ) );
  NAND2_X2 U3375 ( .A1(n4189), .A2(n4188), .ZN(n4187) );
  INV_X2 U3383 ( .A(n3759), .ZN(n4188) );
  NAND2_X2 U3384 ( .A1(n1223), .A2(n347), .ZN(n608) );
  NAND2_X2 U3385 ( .A1(n3451), .A2(n3437), .ZN(n1921) );
  XNOR2_X2 U3387 ( .A(n3424), .B(n3423), .ZN(n3451) );
  NAND2_X2 U3388 ( .A1(n4191), .A2(n4190), .ZN(n2092) );
  NAND2_X2 U3404 ( .A1(n1922), .A2(n3781), .ZN(n4190) );
  NAND2_X2 U3417 ( .A1(n1924), .A2(n1925), .ZN(n4191) );
  NAND2_X2 U3418 ( .A1(n3431), .A2(n100), .ZN(n3411) );
  NOR2_X2 U3419 ( .A1(n3494), .A2(n3760), .ZN(n511) );
  NAND2_X2 U3421 ( .A1(n513), .A2(n512), .ZN(n3494) );
  NAND2_X2 U3427 ( .A1(n2029), .A2(n3232), .ZN(n3231) );
  NAND2_X2 U3428 ( .A1(n1037), .A2(n4192), .ZN(n2029) );
  OAI22_X2 U3432 ( .A1(n3026), .A2(n2828), .B1(n2827), .B2(n2049), .ZN(n710)
         );
  NAND3_X2 U3441 ( .A1(n1036), .A2(n644), .A3(n3226), .ZN(n4192) );
  AND2_X4 U3456 ( .A1(b[1]), .A2(n3176), .ZN(n2384) );
  NOR2_X2 U3458 ( .A1(n4193), .A2(n2279), .ZN(n163) );
  INV_X2 U3484 ( .A(n675), .ZN(n4193) );
  AOI22_X2 U3489 ( .A1(n362), .A2(n363), .B1(n360), .B2(n2128), .ZN(n675) );
  NAND3_X2 U3492 ( .A1(n2072), .A2(n2855), .A3(n2362), .ZN(n1681) );
  NAND3_X2 U3493 ( .A1(n1891), .A2(n1888), .A3(n2360), .ZN(n2072) );
  NAND2_X2 U3497 ( .A1(n4194), .A2(n2974), .ZN(n564) );
  NAND2_X2 U3512 ( .A1(n2973), .A2(n1683), .ZN(n4194) );
  INV_X2 U3516 ( .A(n4195), .ZN(n720) );
  NAND2_X2 U3520 ( .A1(n1483), .A2(n686), .ZN(n4195) );
  INV_X4 U3531 ( .A(n4196), .ZN(n1697) );
  NAND2_X2 U3537 ( .A1(n411), .A2(n3283), .ZN(n4196) );
  NAND2_X2 U3553 ( .A1(n1841), .A2(n1165), .ZN(n2949) );
  NOR2_X2 U3564 ( .A1(n1182), .A2(n4197), .ZN(n2014) );
  OAI22_X1 U3565 ( .A1(n4198), .A2(n2136), .B1(n2931), .B2(n1287), .ZN(n2933)
         );
  INV_X2 U3567 ( .A(n3181), .ZN(n797) );
  NAND2_X2 U3569 ( .A1(n798), .A2(n799), .ZN(n3181) );
  NOR2_X2 U3577 ( .A1(n527), .A2(n2875), .ZN(n2877) );
  NAND2_X2 U3580 ( .A1(n629), .A2(n630), .ZN(n527) );
  NOR2_X1 U3581 ( .A1(n2983), .A2(a[17]), .ZN(n2) );
  NAND2_X2 U3582 ( .A1(n4200), .A2(n4199), .ZN(n365) );
  INV_X2 U3583 ( .A(n3297), .ZN(n4199) );
  INV_X2 U3588 ( .A(n2146), .ZN(n4200) );
  NAND2_X2 U3603 ( .A1(n4201), .A2(n808), .ZN(n2305) );
  NAND3_X2 U3604 ( .A1(n546), .A2(n547), .A3(n1956), .ZN(n4201) );
  NAND2_X2 U3606 ( .A1(n4202), .A2(n254), .ZN(n1627) );
  INV_X1 U3617 ( .A(n1873), .ZN(n2502) );
  OR2_X2 U3621 ( .A1(n3247), .A2(n1842), .ZN(n4204) );
  OR2_X2 U3630 ( .A1(n2564), .A2(n324), .ZN(n4205) );
  AND2_X2 U3631 ( .A1(n3317), .A2(n3318), .ZN(n4206) );
  INV_X1 U3635 ( .A(n1702), .ZN(n1293) );
  NAND2_X2 U3638 ( .A1(n1346), .A2(n1812), .ZN(n201) );
  OR2_X1 U3660 ( .A1(n3893), .A2(n3897), .ZN(n4207) );
  INV_X2 U3668 ( .A(n1984), .ZN(n1409) );
  INV_X4 U885 ( .A(n3453), .ZN(n1121) );
  NOR2_X2 U2967 ( .A1(n843), .A2(n2616), .ZN(n2722) );
  NOR2_X2 U3102 ( .A1(n3429), .A2(n3428), .ZN(n1750) );
  NAND2_X2 U1332 ( .A1(n1279), .A2(n1278), .ZN(n1396) );
  NAND2_X2 U451 ( .A1(n973), .A2(n972), .ZN(n1809) );
  NAND2_X2 U863 ( .A1(n218), .A2(n1565), .ZN(n2967) );
  NAND2_X2 U1213 ( .A1(n375), .A2(n51), .ZN(n1984) );
  NOR2_X1 U51 ( .A1(n2518), .A2(n2517), .ZN(n2202) );
  NAND2_X1 U72 ( .A1(n2384), .A2(n2697), .ZN(n1879) );
  INV_X2 U99 ( .A(n2219), .ZN(n1166) );
  NAND2_X1 U100 ( .A1(n1121), .A2(n56), .ZN(n911) );
  NAND2_X1 U271 ( .A1(n3034), .A2(n55), .ZN(n2076) );
  XOR2_X1 U277 ( .A(n94), .B(n3498), .Z(n440) );
  AND2_X2 U289 ( .A1(n1659), .A2(a[17]), .ZN(n438) );
  BUF_X2 U317 ( .A(n3389), .Z(n1652) );
  NAND2_X1 U368 ( .A1(n2980), .A2(n1554), .ZN(n204) );
  MUX2_X1 U457 ( .A(a[25]), .B(n2145), .S(n3065), .Z(n2570) );
  NAND2_X1 U458 ( .A1(n50), .A2(n4033), .ZN(n1932) );
  INV_X1 U606 ( .A(n358), .ZN(n769) );
  INV_X1 U628 ( .A(n2473), .ZN(n2472) );
  INV_X2 U684 ( .A(n1809), .ZN(n1564) );
  NAND2_X1 U740 ( .A1(n1209), .A2(n56), .ZN(n569) );
  AOI22_X1 U755 ( .A1(n189), .A2(n2563), .B1(n2562), .B2(n69), .ZN(n2526) );
  NAND2_X1 U881 ( .A1(n99), .A2(n3200), .ZN(n1971) );
  INV_X2 U1151 ( .A(n2630), .ZN(n1432) );
  NAND2_X1 U1191 ( .A1(n2064), .A2(n2771), .ZN(n840) );
  NAND2_X1 U1280 ( .A1(n2683), .A2(n2682), .ZN(n2734) );
  NAND2_X1 U1281 ( .A1(n33), .A2(n32), .ZN(n3072) );
  INV_X1 U1670 ( .A(n926), .ZN(n595) );
  INV_X2 U1683 ( .A(n1329), .ZN(n398) );
  NAND2_X1 U1792 ( .A1(n90), .A2(n1649), .ZN(n517) );
  INV_X2 U1802 ( .A(n2262), .ZN(n829) );
  NAND2_X1 U1806 ( .A1(n2602), .A2(n2250), .ZN(n480) );
  NAND3_X1 U1869 ( .A1(n3752), .A2(n3754), .A3(n890), .ZN(n889) );
  INV_X1 U1915 ( .A(n3484), .ZN(n3485) );
  OR2_X1 U2035 ( .A1(n3450), .A2(n3449), .ZN(n3437) );
  OAI21_X1 U2124 ( .B1(n3481), .B2(n3494), .A(n1966), .ZN(n1965) );
  NAND2_X1 U2368 ( .A1(n1495), .A2(n3820), .ZN(n3821) );
  INV_X1 U2439 ( .A(n2748), .ZN(n2749) );
  NOR2_X1 U2532 ( .A1(n2725), .A2(n2724), .ZN(n2748) );
  AND2_X2 U2692 ( .A1(n2758), .A2(n2757), .ZN(n4208) );
  OR2_X1 U2719 ( .A1(n3340), .A2(n3042), .ZN(n4209) );
  OR2_X2 U2746 ( .A1(n2500), .A2(n2309), .ZN(n4210) );
  INV_X2 U2790 ( .A(n3803), .ZN(n3805) );
  INV_X8 U402 ( .A(n3392), .ZN(n3306) );
  NOR2_X4 U617 ( .A1(n160), .A2(n159), .ZN(n3352) );
  INV_X1 U2510 ( .A(n4010), .ZN(n4005) );
  INV_X1 U1752 ( .A(n59), .ZN(n1479) );
  INV_X2 U15 ( .A(n4211), .ZN(n1525) );
  NOR2_X2 U19 ( .A1(n3980), .A2(n3979), .ZN(n4211) );
  INV_X1 U34 ( .A(n3826), .ZN(n3831) );
  NAND2_X1 U35 ( .A1(n59), .A2(n1502), .ZN(n3826) );
  INV_X1 U52 ( .A(n3959), .ZN(n4212) );
  NOR2_X2 U103 ( .A1(n4212), .A2(n3960), .ZN(n282) );
  INV_X1 U109 ( .A(n4021), .ZN(n4213) );
  NOR2_X2 U126 ( .A1(n4213), .A2(n3629), .ZN(n2398) );
  OR2_X2 U172 ( .A1(n4011), .A2(n4009), .ZN(n4013) );
  AND2_X2 U184 ( .A1(n1620), .A2(n1447), .ZN(n3945) );
  AND3_X1 U197 ( .A1(n4010), .A2(n1202), .A3(n1892), .ZN(n3986) );
  OR2_X2 U203 ( .A1(n1350), .A2(n1657), .ZN(n3780) );
  INV_X1 U205 ( .A(n296), .ZN(n3827) );
  NAND2_X1 U209 ( .A1(n3793), .A2(n3792), .ZN(n296) );
  OR2_X2 U213 ( .A1(n3884), .A2(n3825), .ZN(n3888) );
  OAI21_X1 U214 ( .B1(n3840), .B2(n3842), .A(n4214), .ZN(n3850) );
  AOI22_X1 U216 ( .A1(n3843), .A2(n3844), .B1(n3840), .B2(n4215), .ZN(n4214)
         );
  INV_X1 U231 ( .A(n3841), .ZN(n4215) );
  AND2_X2 U234 ( .A1(n68), .A2(n3093), .ZN(n1392) );
  INV_X1 U236 ( .A(n4150), .ZN(n4216) );
  NOR2_X2 U237 ( .A1(n3567), .A2(n4216), .ZN(n4032) );
  AND2_X2 U250 ( .A1(n3646), .A2(n3639), .ZN(n3840) );
  OR2_X2 U305 ( .A1(n3086), .A2(n65), .ZN(n1004) );
  AOI21_X1 U328 ( .B1(n2296), .B2(n3589), .A(n4217), .ZN(n3646) );
  OAI22_X1 U330 ( .A1(n3589), .A2(n4218), .B1(n3643), .B2(n1705), .ZN(n4217)
         );
  INV_X1 U331 ( .A(n2654), .ZN(n4218) );
  AND2_X2 U345 ( .A1(n3439), .A2(n3444), .ZN(n1922) );
  INV_X1 U351 ( .A(n3482), .ZN(n3483) );
  NOR2_X1 U354 ( .A1(n3484), .A2(n3486), .ZN(n3482) );
  AND2_X2 U355 ( .A1(n1383), .A2(n3443), .ZN(n3439) );
  INV_X2 U359 ( .A(n4219), .ZN(n841) );
  NOR2_X2 U364 ( .A1(n2064), .A2(n2771), .ZN(n4219) );
  INV_X2 U377 ( .A(n4220), .ZN(n4147) );
  NOR2_X2 U380 ( .A1(n598), .A2(n3397), .ZN(n4220) );
  INV_X1 U394 ( .A(n4221), .ZN(n1470) );
  NOR2_X2 U396 ( .A1(n1874), .A2(n201), .ZN(n4221) );
  OR2_X2 U425 ( .A1(n3450), .A2(n3449), .ZN(n1546) );
  INV_X2 U462 ( .A(n4222), .ZN(n1127) );
  NOR2_X2 U472 ( .A1(n1382), .A2(n1298), .ZN(n4222) );
  OR2_X2 U525 ( .A1(n2510), .A2(n2509), .ZN(n2422) );
  OAI21_X1 U529 ( .B1(n205), .B2(n3513), .A(n4223), .ZN(n3479) );
  AOI22_X1 U743 ( .A1(n58), .A2(n1088), .B1(n205), .B2(n4224), .ZN(n4223) );
  INV_X1 U800 ( .A(n3512), .ZN(n4224) );
  OR2_X2 U810 ( .A1(n3466), .A2(n3465), .ZN(n3462) );
  AND2_X2 U946 ( .A1(n2429), .A2(n2428), .ZN(n2488) );
  INV_X2 U987 ( .A(n4225), .ZN(n4165) );
  NOR2_X2 U988 ( .A1(n619), .A2(n2961), .ZN(n4225) );
  OAI21_X1 U1019 ( .B1(n90), .B2(n923), .A(n4226), .ZN(n3320) );
  NAND2_X1 U1053 ( .A1(n3430), .A2(n90), .ZN(n4226) );
  OR2_X2 U1078 ( .A1(n2579), .A2(n53), .ZN(n1491) );
  OR2_X2 U1126 ( .A1(n2620), .A2(n2619), .ZN(n2622) );
  OAI21_X1 U1357 ( .B1(n2900), .B2(n2899), .A(n4227), .ZN(n439) );
  INV_X1 U1360 ( .A(n2989), .ZN(n4227) );
  AOI22_X1 U1373 ( .A1(n2902), .A2(n2997), .B1(n3010), .B2(n2901), .ZN(n2989)
         );
  OR2_X2 U1391 ( .A1(n3277), .A2(n1630), .ZN(n1957) );
  INV_X1 U1396 ( .A(n3401), .ZN(n4228) );
  NAND2_X2 U1405 ( .A1(n4228), .A2(n2323), .ZN(n23) );
  INV_X2 U1406 ( .A(n4229), .ZN(n613) );
  OAI211_X1 U1412 ( .C1(n3303), .C2(n205), .A(n1034), .B(n1033), .ZN(n4229) );
  INV_X1 U1417 ( .A(n4230), .ZN(n3390) );
  AOI22_X1 U1420 ( .A1(n1016), .A2(n99), .B1(n1784), .B2(n3472), .ZN(n4230) );
  OAI21_X1 U1429 ( .B1(a[3]), .B2(n3303), .A(n4231), .ZN(n1150) );
  NAND2_X1 U1430 ( .A1(n99), .A2(n1766), .ZN(n4231) );
  NAND2_X2 U1431 ( .A1(n264), .A2(n2507), .ZN(n263) );
  OR2_X2 U1432 ( .A1(n1480), .A2(n2869), .ZN(n1915) );
  INV_X2 U1478 ( .A(n4232), .ZN(n2473) );
  NOR2_X2 U1479 ( .A1(n2469), .A2(n2468), .ZN(n4232) );
  INV_X1 U1480 ( .A(n4233), .ZN(n2495) );
  AOI22_X1 U1483 ( .A1(a[21]), .A2(n3323), .B1(n3217), .B2(n3329), .ZN(n4233)
         );
  OR2_X2 U1484 ( .A1(n2758), .A2(n2757), .ZN(n1251) );
  INV_X2 U1493 ( .A(n4234), .ZN(n842) );
  NOR2_X2 U1499 ( .A1(n2612), .A2(n2611), .ZN(n4234) );
  INV_X1 U1510 ( .A(n725), .ZN(n2517) );
  AOI22_X1 U1511 ( .A1(a[21]), .A2(n3454), .B1(n3455), .B2(n3217), .ZN(n725)
         );
  INV_X1 U1512 ( .A(n4235), .ZN(n2302) );
  AOI22_X1 U1541 ( .A1(n54), .A2(n1237), .B1(n97), .B2(n2084), .ZN(n4235) );
  INV_X2 U1544 ( .A(n4236), .ZN(n2720) );
  AOI22_X1 U1546 ( .A1(a[21]), .A2(n2022), .B1(n3217), .B2(n2980), .ZN(n4236)
         );
  AOI22_X1 U1552 ( .A1(n3109), .A2(n3329), .B1(a[20]), .B2(n3323), .ZN(n460)
         );
  AOI22_X1 U1555 ( .A1(n3128), .A2(n2296), .B1(n55), .B2(n2654), .ZN(n4048) );
  OR2_X2 U1570 ( .A1(n2887), .A2(n1751), .ZN(n632) );
  OR2_X2 U1582 ( .A1(n1751), .A2(n2886), .ZN(n2131) );
  INV_X2 U1583 ( .A(n4237), .ZN(n2616) );
  AOI22_X1 U1584 ( .A1(a[24]), .A2(n1261), .B1(n3589), .B2(n85), .ZN(n4237) );
  INV_X1 U1585 ( .A(n4238), .ZN(n2360) );
  AOI22_X1 U1607 ( .A1(a[14]), .A2(n4075), .B1(n1928), .B2(n2438), .ZN(n4238)
         );
  AOI22_X1 U1609 ( .A1(n98), .A2(n2654), .B1(n2407), .B2(n2296), .ZN(n355) );
  OAI22_X1 U1610 ( .A1(n3475), .A2(n3328), .B1(n58), .B2(n2084), .ZN(n495) );
  INV_X2 U1624 ( .A(n4239), .ZN(n3309) );
  AOI22_X1 U1633 ( .A1(n2045), .A2(n2354), .B1(a[1]), .B2(n86), .ZN(n4239) );
  OR2_X2 U1663 ( .A1(n3216), .A2(n3215), .ZN(n3260) );
  INV_X2 U1681 ( .A(n4240), .ZN(n1949) );
  OAI22_X1 U1682 ( .A1(n3311), .A2(n37), .B1(n3310), .B2(n2057), .ZN(n4240) );
  INV_X1 U1691 ( .A(n4241), .ZN(n1819) );
  AOI22_X1 U1707 ( .A1(n3109), .A2(n3455), .B1(n3454), .B2(a[20]), .ZN(n4241)
         );
  NAND3_X1 U1720 ( .A1(n2145), .A2(n2506), .A3(n1245), .ZN(n2807) );
  INV_X1 U1721 ( .A(n2333), .ZN(n1245) );
  AND2_X2 U1754 ( .A1(n2221), .A2(n2222), .ZN(n2220) );
  OR2_X2 U1755 ( .A1(n3008), .A2(a[14]), .ZN(n4088) );
  INV_X1 U1757 ( .A(n4242), .ZN(n2435) );
  AOI22_X1 U1765 ( .A1(n1554), .A2(n3328), .B1(a[17]), .B2(n2084), .ZN(n4242)
         );
  AOI21_X1 U1775 ( .B1(n1231), .B2(n3124), .A(n4244), .ZN(n2311) );
  NOR2_X1 U1778 ( .A1(n3203), .A2(n1554), .ZN(n4244) );
  OAI22_X1 U1843 ( .A1(n2332), .A2(a[17]), .B1(n2335), .B2(n1554), .ZN(n4050)
         );
  AND2_X2 U1848 ( .A1(n2798), .A2(n2802), .ZN(n2800) );
  OR2_X2 U1855 ( .A1(n3329), .A2(n94), .ZN(n983) );
  OR2_X2 U1886 ( .A1(n3211), .A2(n3306), .ZN(n2213) );
  OR2_X2 U1939 ( .A1(n3016), .A2(n4149), .ZN(n2123) );
  INV_X4 U1960 ( .A(n4245), .ZN(n3709) );
  NAND2_X2 U2025 ( .A1(n3573), .A2(n3574), .ZN(n4245) );
endmodule



    module conf_int_mul__noFF__arch_agnos__w_wrapper_OP_BITWIDTH18_DATA_PATH_BITWIDTH26__acc ( 
        A_in_to_wrapper, B_in_to_wrapper, state_in_to_wrapper, rstP, clk, racc, 
        rapx, P, count0, state_out_of_wrapper, d_internal__apx, acc__sel, 
        A_out, B_out);
  input [25:0] A_in_to_wrapper;
  input [14:0] B_in_to_wrapper;
  input [2:0] state_in_to_wrapper;
  output [31:0] P;
  input [8:0] count0;
  output [2:0] state_out_of_wrapper;
  input [24:0] d_internal__apx;
  output [25:0] A_out;
  output [14:0] B_out;
  //output [24:0] A_out_proc;
  input rstP, clk, racc, rapx, acc__sel;
  wire   n477, n489, n204, n443, n218, n388, n412, n237, n462, n505, n234,
         n464, n235, n451, n233, n478, n244, n449, n501, n214, n406, n229,
         n453, n509, n228, n457, n510, n232, n455, n508, n238, n427, n231,
         n425, n399, net23470, n461, n400, n454, N109, N101, n452, n145, n450,
         n447, n379, n459, n458, n481, N92, n143, n442, N93, N95, N96, n226,
         n335, N97, N111, n465, n230, n435, n217, n467, n391, n227, n460, n511,
         n147, n240, n429, n236, n436, n221, n431, n222, n336, n207, n434,
         n220, n499, n243, n430, n216, n403, n212, n392, n241, n426, n209,
         n423, n223, n338, n239, n428, n208, n439, n215, n398, n225, n433,
         n397, n224, n432, n213, n469, n219, n446, n210, n438, n211, n476,
         n205, n437, n242, n466, d_internal__acc_16, d_internal__acc_13, n417,
         d_internal__acc_10, d_internal__acc_14, d_internal__acc_11,
         d_internal__acc_9, d_internal__acc_8, n255, n256, d_internal__acc_12,
         n401, d_internal__acc_17, n421, n271, n18, n164, n419, n479, n424,
         n488, n487, n486, n483, n484, n474, n480, n471, n448, n473, n445,
         n456, d_internal__acc_18, n196, n206, n270, n120, n121, n122, n124,
         n128, n129, n131, n133, n134, n136, n138, n139, n482, n141, n142,
         n144, n485, n148, n149, n150, n151, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n197, n198,
         n199, n200, n201, n202, n203, n245, n246, n247, n248, n249, n250,
         n251, n253, n254, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n272, n273, n274, n275, n276, n277,
         n278, n281, n282, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n337, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n380, n381, n382, n383, n384, n385,
         n386, n387, n389, n390, n393, n394, n395, n396, n404, n405, n407,
         n408, n409, n410, n411, n413, n414, n415, n416, n418, n420, n422,
         n440, n441, n444, n463, n468, n470, n472, n490;
  wire   [39:20] d_internal__acc;
  //assign A_out_proc[22] = n445;

  DFFR_X2 \b_reg_reg[0]  ( .D(n204), .CK(clk), .RN(n422), .QN(n443), .Q() );
  DFFR_X2 \b_reg_reg[14]  ( .D(n218), .CK(clk), .RN(n468), .QN(n388), .Q(n412)
         );
  DFFR_X2 \a_reg_reg[18]  ( .D(n237), .CK(clk), .RN(n440), .QN(n462), .Q(n505)
         );
  DFFR_X2 \a_reg_reg[15]  ( .D(n234), .CK(clk), .RN(n440), .QN(n464), .Q(
        A_out[15]) );
  DFFR_X2 \a_reg_reg[16]  ( .D(n235), .CK(clk), .RN(n463), .QN(n451), .Q(
        A_out[16]) );
  DFFR_X2 \a_reg_reg[14]  ( .D(n233), .CK(clk), .RN(n440), .QN(n478), .Q(
        A_out[14]) );
  DFFR_X2 \a_reg_reg[25]  ( .D(n244), .CK(clk), .RN(n420), .QN(n449), .Q(n501)
         );
  DFFR_X2 \b_reg_reg[10]  ( .D(n214), .CK(clk), .RN(n418), .QN(n406), .Q(
        B_out[10]) );
  DFFR_X2 \a_reg_reg[10]  ( .D(n229), .CK(clk), .RN(n422), .QN(n453), .Q(n509)
         );
  DFFR_X2 \a_reg_reg[9]  ( .D(n228), .CK(clk), .RN(n422), .QN(n457), .Q(n510)
         );
  DFFR_X2 \a_reg_reg[13]  ( .D(n232), .CK(clk), .RN(n444), .QN(n455), .Q(n508)
         );
  DFFR_X2 \a_reg_reg[19]  ( .D(n238), .CK(clk), .RN(n422), .QN(n427), .Q(
        A_out[19]) );
  DFFR_X2 \a_reg_reg[12]  ( .D(n231), .CK(clk), .RN(n444), .QN(n425), .Q(
        A_out[12]) );
  DFFR_X1 \c_reg_reg[4]  ( .D(n399), .CK(clk), .RN(net23470), .QN(), .Q(P[4])
         );
  DFFR_X1 \c_reg_reg[16]  ( .D(n461), .CK(clk), .RN(net23470), .QN(), .Q(P[16]) );
  DFFR_X1 \c_reg_reg[20]  ( .D(n470), .CK(clk), .RN(net23470), .QN(), .Q(P[20]) );
  DFFR_X1 \c_reg_reg[31]  ( .D(n400), .CK(clk), .RN(net23470), .QN(), .Q(P[31]) );
  DFFR_X1 \c_reg_reg[21]  ( .D(n454), .CK(clk), .RN(net23470), .QN(), .Q(P[21]) );
  DFFR_X1 \c_reg_reg[25]  ( .D(N109), .CK(clk), .RN(net23470), .QN(), .Q(P[25]) );
  DFFR_X1 \c_reg_reg[17]  ( .D(N101), .CK(clk), .RN(net23470), .QN(), .Q(P[17]) );
  DFFR_X1 \c_reg_reg[26]  ( .D(n452), .CK(clk), .RN(net23470), .QN(), .Q(P[26]) );
  DFFR_X1 \c_reg_reg[18]  ( .D(n145), .CK(clk), .RN(net23470), .QN(), .Q(P[18]) );
  DFFR_X1 \c_reg_reg[19]  ( .D(n450), .CK(clk), .RN(net23470), .QN(), .Q(P[19]) );
  DFFR_X1 \c_reg_reg[15]  ( .D(n472), .CK(clk), .RN(net23470), .QN(), .Q(P[15]) );
  DFFR_X1 \c_reg_reg[14]  ( .D(n447), .CK(clk), .RN(net23470), .QN(), .Q(P[14]) );
  DFFR_X1 \c_reg_reg[29]  ( .D(n379), .CK(clk), .RN(net23470), .QN(), .Q(P[29]) );
  DFFR_X1 \c_reg_reg[23]  ( .D(n459), .CK(clk), .RN(net23470), .QN(), .Q(P[23]) );
  DFFR_X1 \c_reg_reg[22]  ( .D(n458), .CK(clk), .RN(net23470), .QN(), .Q(P[22]) );
  DFFR_X1 \c_reg_reg[24]  ( .D(n481), .CK(clk), .RN(net23470), .QN(), .Q(P[24]) );
  DFFR_X1 \c_reg_reg[8]  ( .D(N92), .CK(clk), .RN(net23470), .QN(), .Q(P[8])
         );
  DFFR_X1 \c_reg_reg[7]  ( .D(n143), .CK(clk), .RN(net23470), .QN(), .Q(P[7])
         );
  DFFR_X1 \c_reg_reg[10]  ( .D(n442), .CK(clk), .RN(net23470), .QN(), .Q(P[10]) );
  DFFR_X1 \c_reg_reg[9]  ( .D(N93), .CK(clk), .RN(net23470), .QN(), .Q(P[9])
         );
  DFFR_X1 \c_reg_reg[11]  ( .D(N95), .CK(clk), .RN(net23470), .QN(), .Q(P[11])
         );
  DFFR_X1 \c_reg_reg[12]  ( .D(N96), .CK(clk), .RN(net23470), .QN(), .Q(P[12])
         );
  DFFR_X2 \a_reg_reg[7]  ( .D(n226), .CK(clk), .RN(n441), .QN(n335), .Q() );
  DFFR_X1 \c_reg_reg[13]  ( .D(N97), .CK(clk), .RN(net23470), .QN(), .Q(P[13])
         );
  DFFR_X1 \c_reg_reg[27]  ( .D(N111), .CK(clk), .RN(net23470), .QN(), .Q(P[27]) );
  DFFR_X1 \c_reg_reg[30]  ( .D(n465), .CK(clk), .RN(net23470), .QN(), .Q(P[30]) );
  DFFR_X2 \a_reg_reg[11]  ( .D(n230), .CK(clk), .RN(n422), .QN(n435), .Q(
        A_out[11]) );
  DFFR_X1 \c_reg_reg[28]  ( .D(n467), .CK(clk), .RN(net23470), .QN(), .Q(P[28]) );
  DFFR_X1 \c_reg_reg[5]  ( .D(n391), .CK(clk), .RN(net23470), .QN(), .Q(P[5])
         );
  DFFR_X2 \a_reg_reg[8]  ( .D(n227), .CK(clk), .RN(n420), .QN(n460), .Q(n511)
         );
  DFFR_X1 \c_reg_reg[6]  ( .D(n147), .CK(clk), .RN(net23470), .QN(P[6]), .Q()
         );
  DFFR_X2 \a_reg_reg[17]  ( .D(n236), .CK(clk), .RN(n416), .QN(n436), .Q(
        A_out[17]) );
  DFFR_X2 \a_reg_reg[3]  ( .D(n222), .CK(clk), .RN(n420), .QN(n336), .Q() );
  DFFR_X2 \b_reg_reg[3]  ( .D(n207), .CK(clk), .RN(n418), .QN(n434), .Q(
        B_out[3]) );
  DFFR_X2 \a_reg_reg[1]  ( .D(n220), .CK(clk), .RN(n420), .QN(n499), .Q() );
  DFFR_X2 \a_reg_reg[24]  ( .D(n243), .CK(clk), .RN(n441), .QN(n430), .Q(
        A_out[24]) );
  DFFR_X2 \b_reg_reg[12]  ( .D(n216), .CK(clk), .RN(n440), .QN(n403), .Q(
        B_out[12]) );
  DFFR_X2 \b_reg_reg[8]  ( .D(n212), .CK(clk), .RN(n418), .QN(n392), .Q(
        B_out[8]) );
  DFFR_X2 \a_reg_reg[22]  ( .D(n241), .CK(clk), .RN(n468), .QN(n426), .Q(
        A_out[22]) );
  DFFR_X1 \a_reg_reg[4]  ( .D(n223), .CK(clk), .RN(n441), .QN(n338), .Q(
        A_out[4]) );
  DFFR_X2 \a_reg_reg[20]  ( .D(n239), .CK(clk), .RN(n440), .QN(n428), .Q(
        A_out[20]) );
  DFFR_X2 \b_reg_reg[4]  ( .D(n208), .CK(clk), .RN(n416), .QN(n439), .Q(
        B_out[4]) );
  DFFR_X2 \b_reg_reg[11]  ( .D(n215), .CK(clk), .RN(n418), .QN(n398), .Q(
        B_out[11]) );
  DFFR_X1 \a_reg_reg[6]  ( .D(n225), .CK(clk), .RN(n441), .QN(n433), .Q(
        A_out[6]) );
  DFFR_X1 \state_reg[0]  ( .D(state_in_to_wrapper[0]), .CK(clk), .RN(n468), 
        .QN(n397), .Q(state_out_of_wrapper[0]) );
  DFFR_X1 \a_reg_reg[5]  ( .D(n224), .CK(clk), .RN(n463), .QN(n432), .Q(
        A_out[5]) );
  DFFR_X2 \b_reg_reg[9]  ( .D(n213), .CK(clk), .RN(n418), .QN(n469), .Q(
        B_out[9]) );
  DFFR_X1 \a_reg_reg[0]  ( .D(n219), .CK(clk), .RN(n420), .QN(n446), .Q(
        A_out[0]) );
  DFFR_X2 \b_reg_reg[7]  ( .D(n211), .CK(clk), .RN(n416), .QN(n476), .Q(
        B_out[7]) );
  DFFR_X1 \c_reg_reg[2]  ( .D(n270), .CK(clk), .RN(net23470), .QN(P[2]), .Q()
         );
  DFFR_X1 \c_reg_reg[3]  ( .D(n271), .CK(clk), .RN(net23470), .QN(P[3]), .Q()
         );
  DFFR_X2 \b_reg_reg[2]  ( .D(n206), .CK(clk), .RN(n468), .QN(n196), .Q(
        B_out[2]) );
  DFFR_X2 \b_reg_reg[6]  ( .D(n210), .CK(clk), .RN(n416), .QN(n438), .Q(
        B_out[6]) );
  DFFR_X2 \b_reg_reg[5]  ( .D(n209), .CK(clk), .RN(n416), .QN(n423), .Q(
        B_out[5]) );
  DFFR_X1 \state_reg[1]  ( .D(state_in_to_wrapper[1]), .CK(clk), .RN(n463), 
        .QN(), .Q(state_out_of_wrapper[1]) );
  DFFR_X2 \b_reg_reg[1]  ( .D(n205), .CK(clk), .RN(n468), .QN(n437), .Q(
        B_out[1]) );
  DFFR_X2 \b_reg_reg[13]  ( .D(n217), .CK(clk), .RN(n444), .QN(n415), .Q(n477)
         );
  DFFR_X1 \a_reg_reg[21]  ( .D(n240), .CK(clk), .RN(n441), .QN(n429), .Q(
        A_out[21]) );
  DFFR_X1 \state_reg[2]  ( .D(state_in_to_wrapper[2]), .CK(clk), .RN(n463), 
        .QN(), .Q(state_out_of_wrapper[2]) );
  DFFR_X1 \a_reg_reg[23]  ( .D(n242), .CK(clk), .RN(n444), .QN(n466), .Q(
        A_out[23]) );
  NAND2_X1 U239 ( .A1(n350), .A2(n327), .ZN(n377) );
  NAND2_X1 U243 ( .A1(n284), .A2(acc__sel), .ZN(n282) );
  NAND2_X1 U245 ( .A1(n351), .A2(n327), .ZN(n376) );
  AOI21_X1 U246 ( .B1(d_internal__acc_18), .B2(n171), .A(n263), .ZN(n268) );
  INV_X1 U247 ( .A(n330), .ZN(n386) );
  INV_X1 U248 ( .A(racc), .ZN(n463) );
  INV_X4 U250 ( .A(n390), .ZN(n350) );
  INV_X8 U252 ( .A(n409), .ZN(n171) );
  INV_X2 U253 ( .A(n282), .ZN(n281) );
  OR2_X2 U256 ( .A1(d_internal__acc[20]), .A2(n414), .ZN(n195) );
  NAND2_X1 U257 ( .A1(n364), .A2(n363), .ZN(N95) );
  INV_X2 U258 ( .A(d_internal__acc_12), .ZN(n292) );
  INV_X2 U259 ( .A(d_internal__acc_16), .ZN(n394) );
  NOR2_X1 U260 ( .A1(n180), .A2(n179), .ZN(n363) );
  AOI22_X1 U261 ( .A1(n266), .A2(n171), .B1(d_internal__apx[4]), .B2(n410), 
        .ZN(n265) );
  AOI22_X1 U262 ( .A1(n359), .A2(n171), .B1(n410), .B2(d_internal__apx[2]), 
        .ZN(n360) );
  INV_X2 U263 ( .A(n417), .ZN(n266) );
  INV_X2 U266 ( .A(d_internal__acc_9), .ZN(n358) );
  AOI22_X1 U269 ( .A1(n411), .A2(d_internal__apx[1]), .B1(n410), .B2(
        d_internal__apx[6]), .ZN(n296) );
  INV_X1 U271 ( .A(n171), .ZN(n181) );
  INV_X1 U272 ( .A(n414), .ZN(n172) );
  AND2_X1 U273 ( .A1(n410), .A2(d_internal__apx[3]), .ZN(n179) );
  NAND2_X1 U275 ( .A1(n410), .A2(d_internal__apx[0]), .ZN(n197) );
  NOR2_X2 U276 ( .A1(n285), .A2(n286), .ZN(n411) );
  NOR2_X2 U277 ( .A1(n315), .A2(n286), .ZN(n410) );
  NOR2_X2 U279 ( .A1(state_out_of_wrapper[2]), .A2(n318), .ZN(n315) );
  INV_X4 U281 ( .A(n478), .ZN(n122) );
  NAND2_X2 U282 ( .A1(state_out_of_wrapper[1]), .A2(n397), .ZN(n318) );
  INV_X4 U283 ( .A(n435), .ZN(n131) );
  INV_X4 U284 ( .A(n436), .ZN(n134) );
  INV_X2 U285 ( .A(n464), .ZN(n120) );
  INV_X2 U286 ( .A(n451), .ZN(n121) );
  INV_X2 U287 ( .A(n462), .ZN(A_out[18]) );
  INV_X2 U288 ( .A(n455), .ZN(A_out[13]) );
  INV_X8 U290 ( .A(n398), .ZN(n148) );
  NAND2_X2 U291 ( .A1(n174), .A2(n173), .ZN(n400) );
  NAND2_X2 U292 ( .A1(d_internal__acc[34]), .A2(n171), .ZN(n173) );
  AOI21_X2 U293 ( .B1(d_internal__acc[39]), .B2(n407), .A(n186), .ZN(n174) );
  NAND2_X2 U295 ( .A1(n201), .A2(n202), .ZN(n452) );
  INV_X4 U296 ( .A(n407), .ZN(n414) );
  NAND2_X2 U297 ( .A1(n315), .A2(n281), .ZN(n409) );
  NOR2_X4 U298 ( .A1(n315), .A2(n282), .ZN(n407) );
  NAND3_X2 U299 ( .A1(n177), .A2(n176), .A3(n395), .ZN(N97) );
  NAND2_X2 U300 ( .A1(n394), .A2(n171), .ZN(n176) );
  NAND2_X2 U301 ( .A1(n178), .A2(n172), .ZN(n177) );
  INV_X2 U302 ( .A(d_internal__acc[21]), .ZN(n178) );
  INV_X2 U303 ( .A(d_internal__acc_14), .ZN(n362) );
  NOR2_X2 U304 ( .A1(d_internal__acc_14), .A2(n181), .ZN(n180) );
  AOI21_X2 U305 ( .B1(n182), .B2(n171), .A(n273), .ZN(n190) );
  INV_X2 U306 ( .A(d_internal__acc[22]), .ZN(n182) );
  NAND2_X2 U307 ( .A1(n183), .A2(n189), .ZN(n458) );
  NAND2_X2 U308 ( .A1(n184), .A2(n172), .ZN(n183) );
  NAND2_X2 U310 ( .A1(d_internal__acc_17), .A2(n171), .ZN(n298) );
  NAND3_X2 U311 ( .A1(n298), .A2(n297), .A3(n296), .ZN(n447) );
  NAND2_X2 U312 ( .A1(n185), .A2(n290), .ZN(N111) );
  NOR2_X2 U313 ( .A1(n289), .A2(n288), .ZN(n185) );
  INV_X2 U314 ( .A(n366), .ZN(n186) );
  NAND2_X2 U315 ( .A1(n188), .A2(n187), .ZN(n470) );
  NAND2_X2 U316 ( .A1(d_internal__acc[28]), .A2(n407), .ZN(n187) );
  AOI21_X2 U317 ( .B1(d_internal__acc[23]), .B2(n171), .A(n203), .ZN(n188) );
  AOI21_X2 U318 ( .B1(d_internal__acc[25]), .B2(n171), .A(n302), .ZN(n189) );
  NAND2_X2 U319 ( .A1(d_internal__acc_17), .A2(n407), .ZN(n294) );
  OAI21_X2 U320 ( .B1(d_internal__acc[27]), .B2(n414), .A(n190), .ZN(n450) );
  OAI21_X2 U321 ( .B1(d_internal__acc[27]), .B2(n409), .A(n191), .ZN(n481) );
  AOI21_X2 U322 ( .B1(d_internal__acc[32]), .B2(n407), .A(n300), .ZN(n191) );
  NAND2_X2 U323 ( .A1(n193), .A2(n192), .ZN(n465) );
  AOI21_X2 U324 ( .B1(d_internal__acc[33]), .B2(n171), .A(n312), .ZN(n192) );
  NAND2_X2 U325 ( .A1(n194), .A2(n407), .ZN(n193) );
  INV_X2 U326 ( .A(d_internal__acc[38]), .ZN(n194) );
  INV_X1 U327 ( .A(n315), .ZN(n285) );
  NAND2_X1 U328 ( .A1(count0[2]), .A2(count0[3]), .ZN(n314) );
  INV_X1 U331 ( .A(n413), .ZN(n261) );
  NAND2_X1 U332 ( .A1(n358), .A2(n407), .ZN(n256) );
  NAND2_X1 U333 ( .A1(d_internal__acc_11), .A2(n407), .ZN(n271) );
  AOI22_X1 U334 ( .A1(n330), .A2(B_out[4]), .B1(n328), .B2(B_in_to_wrapper[4]), 
        .ZN(n329) );
  INV_X1 U335 ( .A(n377), .ZN(n328) );
  OAI21_X1 U336 ( .B1(n175), .B2(n386), .A(n325), .ZN(n212) );
  AOI22_X1 U337 ( .A1(n362), .A2(n407), .B1(n171), .B2(n358), .ZN(n147) );
  NOR2_X1 U338 ( .A1(d_internal__acc_13), .A2(n414), .ZN(n391) );
  INV_X1 U339 ( .A(n408), .ZN(n278) );
  INV_X1 U340 ( .A(n311), .ZN(n312) );
  OAI22_X1 U341 ( .A1(n417), .A2(n414), .B1(d_internal__acc_10), .B2(n409), 
        .ZN(n143) );
  INV_X1 U342 ( .A(n299), .ZN(n300) );
  INV_X1 U343 ( .A(n303), .ZN(n277) );
  INV_X1 U344 ( .A(n365), .ZN(n263) );
  INV_X1 U345 ( .A(n304), .ZN(n305) );
  INV_X1 U346 ( .A(n291), .ZN(n264) );
  INV_X1 U347 ( .A(n309), .ZN(n310) );
  INV_X1 U348 ( .A(n367), .ZN(n259) );
  INV_X1 U349 ( .A(n405), .ZN(n276) );
  INV_X1 U350 ( .A(n295), .ZN(n203) );
  INV_X1 U351 ( .A(n396), .ZN(n275) );
  NOR2_X1 U352 ( .A1(d_internal__acc_12), .A2(n414), .ZN(n399) );
  INV_X4 U353 ( .A(n335), .ZN(A_out[7]) );
  INV_X4 U354 ( .A(n457), .ZN(A_out[9]) );
  NAND3_X2 U355 ( .A1(n199), .A2(n198), .A3(n197), .ZN(N92) );
  NAND2_X2 U357 ( .A1(n394), .A2(n407), .ZN(n199) );
  OAI21_X2 U358 ( .B1(d_internal__acc[24]), .B2(n409), .A(n200), .ZN(n454) );
  AOI21_X2 U359 ( .B1(d_internal__acc[29]), .B2(n407), .A(n276), .ZN(n200) );
  NAND2_X2 U360 ( .A1(d_internal__acc[34]), .A2(n407), .ZN(n201) );
  AOI21_X1 U361 ( .B1(d_internal__acc[29]), .B2(n171), .A(n264), .ZN(n202) );
  NAND2_X2 U362 ( .A1(n246), .A2(n245), .ZN(N109) );
  NAND2_X2 U363 ( .A1(d_internal__acc[28]), .A2(n171), .ZN(n245) );
  AOI21_X2 U364 ( .B1(d_internal__acc[33]), .B2(n407), .A(n259), .ZN(n246) );
  NAND2_X1 U365 ( .A1(d_internal__acc_18), .A2(n407), .ZN(n361) );
  INV_X1 U366 ( .A(B_out[12]), .ZN(n247) );
  INV_X1 U368 ( .A(B_out[3]), .ZN(n248) );
  NAND2_X1 U369 ( .A1(n407), .A2(d_internal__acc[25]), .ZN(n254) );
  NAND2_X1 U370 ( .A1(n407), .A2(d_internal__acc[26]), .ZN(n307) );
  INV_X4 U371 ( .A(n392), .ZN(n482) );
  OAI21_X1 U372 ( .B1(n249), .B2(n386), .A(n323), .ZN(n215) );
  INV_X4 U373 ( .A(n469), .ZN(n149) );
  OAI21_X2 U374 ( .B1(d_internal__acc[31]), .B2(n414), .A(n272), .ZN(n459) );
  INV_X8 U375 ( .A(n336), .ZN(A_out[3]) );
  INV_X1 U376 ( .A(B_out[11]), .ZN(n249) );
  OAI21_X2 U377 ( .B1(d_internal__acc[31]), .B2(n409), .A(n267), .ZN(n467) );
  INV_X1 U378 ( .A(B_out[7]), .ZN(n250) );
  INV_X1 U379 ( .A(n124), .ZN(n251) );
  INV_X4 U380 ( .A(n415), .ZN(B_out[13]) );
  INV_X1 U381 ( .A(B_out[9]), .ZN(n253) );
  INV_X8 U382 ( .A(n476), .ZN(n150) );
  NAND2_X1 U383 ( .A1(n410), .A2(d_internal__apx[1]), .ZN(n293) );
  AOI22_X1 U384 ( .A1(n411), .A2(d_internal__apx[18]), .B1(n410), .B2(
        d_internal__apx[23]), .ZN(n366) );
  AOI22_X1 U385 ( .A1(n411), .A2(d_internal__apx[7]), .B1(n410), .B2(
        d_internal__apx[12]), .ZN(n295) );
  AOI22_X1 U386 ( .A1(n411), .A2(d_internal__apx[0]), .B1(n410), .B2(
        d_internal__apx[5]), .ZN(n395) );
  AOI22_X1 U387 ( .A1(n411), .A2(d_internal__apx[4]), .B1(n410), .B2(
        d_internal__apx[9]), .ZN(n309) );
  AOI22_X1 U388 ( .A1(n411), .A2(d_internal__apx[5]), .B1(n410), .B2(
        d_internal__apx[10]), .ZN(n304) );
  AOI22_X1 U389 ( .A1(n411), .A2(d_internal__apx[14]), .B1(n410), .B2(
        d_internal__apx[19]), .ZN(n287) );
  AOI22_X1 U390 ( .A1(n411), .A2(d_internal__apx[12]), .B1(n410), .B2(
        d_internal__apx[17]), .ZN(n367) );
  AOI22_X1 U391 ( .A1(n411), .A2(d_internal__apx[17]), .B1(n410), .B2(
        d_internal__apx[22]), .ZN(n311) );
  AOI22_X1 U392 ( .A1(n411), .A2(d_internal__apx[10]), .B1(d_internal__apx[15]), .B2(n410), .ZN(n303) );
  AOI22_X1 U393 ( .A1(n411), .A2(d_internal__apx[2]), .B1(n410), .B2(
        d_internal__apx[7]), .ZN(n365) );
  AOI22_X1 U394 ( .A1(n411), .A2(d_internal__apx[6]), .B1(n410), .B2(
        d_internal__apx[11]), .ZN(n404) );
  AOI22_X1 U395 ( .A1(n411), .A2(d_internal__apx[13]), .B1(n410), .B2(
        d_internal__apx[18]), .ZN(n291) );
  AOI22_X1 U396 ( .A1(n411), .A2(d_internal__apx[16]), .B1(n410), .B2(
        d_internal__apx[21]), .ZN(n413) );
  AOI22_X1 U397 ( .A1(n411), .A2(d_internal__apx[3]), .B1(n410), .B2(
        d_internal__apx[8]), .ZN(n396) );
  AOI22_X1 U398 ( .A1(n411), .A2(d_internal__apx[9]), .B1(n410), .B2(
        d_internal__apx[14]), .ZN(n301) );
  AOI22_X1 U399 ( .A1(n411), .A2(d_internal__apx[15]), .B1(n410), .B2(
        d_internal__apx[20]), .ZN(n408) );
  AOI22_X1 U400 ( .A1(n411), .A2(d_internal__apx[8]), .B1(n410), .B2(
        d_internal__apx[13]), .ZN(n405) );
  AOI22_X1 U401 ( .A1(n411), .A2(d_internal__apx[11]), .B1(n410), .B2(
        d_internal__apx[16]), .ZN(n299) );
  AOI22_X1 U402 ( .A1(n351), .A2(A_in_to_wrapper[0]), .B1(A_in_to_wrapper[8]), 
        .B2(n350), .ZN(n352) );
  AOI22_X1 U403 ( .A1(n351), .A2(B_in_to_wrapper[8]), .B1(B_in_to_wrapper[9]), 
        .B2(n350), .ZN(n349) );
  AOI22_X1 U404 ( .A1(n351), .A2(A_in_to_wrapper[12]), .B1(A_in_to_wrapper[20]), .B2(n350), .ZN(n348) );
  AOI22_X1 U405 ( .A1(n351), .A2(A_in_to_wrapper[14]), .B1(A_in_to_wrapper[22]), .B2(n350), .ZN(n347) );
  AOI22_X1 U406 ( .A1(n351), .A2(A_in_to_wrapper[16]), .B1(A_in_to_wrapper[24]), .B2(n350), .ZN(n346) );
  AOI22_X1 U407 ( .A1(n351), .A2(A_in_to_wrapper[9]), .B1(A_in_to_wrapper[17]), 
        .B2(n350), .ZN(n345) );
  AOI22_X1 U408 ( .A1(n351), .A2(A_in_to_wrapper[13]), .B1(A_in_to_wrapper[21]), .B2(n350), .ZN(n344) );
  AOI22_X1 U409 ( .A1(n351), .A2(A_in_to_wrapper[8]), .B1(A_in_to_wrapper[16]), 
        .B2(n350), .ZN(n343) );
  AOI22_X1 U410 ( .A1(n351), .A2(A_in_to_wrapper[15]), .B1(A_in_to_wrapper[23]), .B2(n350), .ZN(n342) );
  AOI22_X1 U411 ( .A1(n351), .A2(A_in_to_wrapper[5]), .B1(A_in_to_wrapper[13]), 
        .B2(n350), .ZN(n341) );
  AOI22_X1 U412 ( .A1(n351), .A2(A_in_to_wrapper[10]), .B1(A_in_to_wrapper[18]), .B2(n350), .ZN(n340) );
  AOI22_X1 U413 ( .A1(n351), .A2(A_in_to_wrapper[1]), .B1(A_in_to_wrapper[9]), 
        .B2(n350), .ZN(n339) );
  AOI22_X1 U414 ( .A1(n351), .A2(A_in_to_wrapper[17]), .B1(A_in_to_wrapper[25]), .B2(n350), .ZN(n337) );
  AOI22_X1 U415 ( .A1(n351), .A2(A_in_to_wrapper[2]), .B1(A_in_to_wrapper[10]), 
        .B2(n350), .ZN(n334) );
  AOI22_X1 U416 ( .A1(n351), .A2(B_in_to_wrapper[13]), .B1(B_in_to_wrapper[14]), .B2(n350), .ZN(n333) );
  AOI22_X1 U417 ( .A1(n351), .A2(A_in_to_wrapper[11]), .B1(A_in_to_wrapper[19]), .B2(n350), .ZN(n332) );
  AOI22_X1 U418 ( .A1(n351), .A2(B_in_to_wrapper[12]), .B1(B_in_to_wrapper[13]), .B2(n350), .ZN(n331) );
  AOI22_X1 U419 ( .A1(n351), .A2(B_in_to_wrapper[7]), .B1(B_in_to_wrapper[8]), 
        .B2(n350), .ZN(n325) );
  AOI22_X1 U420 ( .A1(n351), .A2(B_in_to_wrapper[10]), .B1(B_in_to_wrapper[11]), .B2(n350), .ZN(n323) );
  AOI22_X1 U421 ( .A1(n351), .A2(B_in_to_wrapper[9]), .B1(B_in_to_wrapper[10]), 
        .B2(n350), .ZN(n326) );
  OAI21_X1 U422 ( .B1(n357), .B2(n415), .A(n331), .ZN(n217) );
  OAI21_X1 U423 ( .B1(n460), .B2(n357), .A(n352), .ZN(n227) );
  OAI21_X1 U424 ( .B1(n253), .B2(n357), .A(n349), .ZN(n213) );
  OAI21_X1 U425 ( .B1(n428), .B2(n357), .A(n348), .ZN(n239) );
  OAI21_X1 U426 ( .B1(n426), .B2(n357), .A(n347), .ZN(n241) );
  OAI21_X1 U427 ( .B1(n430), .B2(n357), .A(n346), .ZN(n243) );
  OAI21_X1 U428 ( .B1(n436), .B2(n357), .A(n345), .ZN(n236) );
  OAI21_X1 U429 ( .B1(n429), .B2(n357), .A(n344), .ZN(n240) );
  OAI21_X1 U430 ( .B1(n451), .B2(n357), .A(n343), .ZN(n235) );
  OAI21_X1 U431 ( .B1(n466), .B2(n357), .A(n342), .ZN(n242) );
  OAI21_X1 U432 ( .B1(n455), .B2(n357), .A(n341), .ZN(n232) );
  OAI21_X1 U433 ( .B1(n462), .B2(n357), .A(n340), .ZN(n237) );
  OAI21_X1 U434 ( .B1(n457), .B2(n357), .A(n339), .ZN(n228) );
  OAI21_X1 U435 ( .B1(n449), .B2(n357), .A(n337), .ZN(n244) );
  OAI21_X1 U436 ( .B1(n453), .B2(n357), .A(n334), .ZN(n229) );
  OAI21_X1 U437 ( .B1(n388), .B2(n357), .A(n333), .ZN(n218) );
  OAI21_X1 U438 ( .B1(n427), .B2(n357), .A(n332), .ZN(n238) );
  OAI22_X1 U439 ( .A1(n357), .A2(n443), .B1(n368), .B2(n377), .ZN(n204) );
  OAI22_X1 U440 ( .A1(n357), .A2(n335), .B1(n377), .B2(n389), .ZN(n226) );
  OAI22_X1 U441 ( .A1(n357), .A2(n446), .B1(n377), .B2(n356), .ZN(n219) );
  OAI22_X1 U442 ( .A1(n357), .A2(n338), .B1(n377), .B2(n382), .ZN(n223) );
  OAI22_X1 U443 ( .A1(n357), .A2(n433), .B1(n377), .B2(n384), .ZN(n225) );
  OAI22_X1 U444 ( .A1(n357), .A2(n499), .B1(n377), .B2(n355), .ZN(n220) );
  OAI22_X1 U445 ( .A1(n357), .A2(n336), .B1(n377), .B2(n380), .ZN(n222) );
  OAI22_X1 U446 ( .A1(n357), .A2(n432), .B1(n377), .B2(n353), .ZN(n224) );
  INV_X4 U447 ( .A(n439), .ZN(n485) );
  NAND2_X2 U448 ( .A1(n257), .A2(n254), .ZN(N101) );
  NOR2_X2 U449 ( .A1(n258), .A2(n310), .ZN(n257) );
  NOR2_X2 U450 ( .A1(d_internal__acc[20]), .A2(n409), .ZN(n258) );
  OAI21_X2 U451 ( .B1(d_internal__acc[37]), .B2(n414), .A(n260), .ZN(n379) );
  AOI21_X2 U452 ( .B1(d_internal__acc[32]), .B2(n171), .A(n261), .ZN(n260) );
  NAND3_X2 U453 ( .A1(n262), .A2(n294), .A3(n293), .ZN(N93) );
  NAND2_X2 U454 ( .A1(n292), .A2(n171), .ZN(n262) );
  NAND2_X2 U455 ( .A1(n265), .A2(n195), .ZN(N96) );
  AOI21_X2 U456 ( .B1(d_internal__acc[36]), .B2(n407), .A(n278), .ZN(n267) );
  NAND2_X2 U457 ( .A1(n269), .A2(n268), .ZN(n472) );
  AOI21_X2 U458 ( .B1(d_internal__acc[26]), .B2(n171), .A(n277), .ZN(n272) );
  OAI21_X2 U459 ( .B1(d_internal__acc[24]), .B2(n414), .A(n274), .ZN(n461) );
  AOI21_X2 U460 ( .B1(n164), .B2(n171), .A(n275), .ZN(n274) );
  //INV_X1 U461 ( .A(n401), .ZN(A_out_proc[23]) );
  OAI21_X1 U462 ( .B1(n376), .B2(n371), .A(n329), .ZN(n208) );
  INV_X1 U463 ( .A(racc), .ZN(n468) );
  INV_X1 U464 ( .A(racc), .ZN(n441) );
  INV_X1 U465 ( .A(racc), .ZN(n420) );
  INV_X1 U466 ( .A(racc), .ZN(n422) );
  INV_X1 U467 ( .A(racc), .ZN(n440) );
  INV_X1 U468 ( .A(racc), .ZN(n416) );
  INV_X1 U469 ( .A(racc), .ZN(n418) );
  INV_X1 U470 ( .A(racc), .ZN(n444) );
  NAND2_X1 U471 ( .A1(state_out_of_wrapper[2]), .A2(state_out_of_wrapper[0]), 
        .ZN(n321) );
  INV_X1 U472 ( .A(B_in_to_wrapper[1]), .ZN(n369) );
  NAND2_X1 U473 ( .A1(n164), .A2(n407), .ZN(n364) );
  INV_X1 U474 ( .A(A_in_to_wrapper[6]), .ZN(n384) );
  OAI22_X1 U475 ( .A1(n357), .A2(n431), .B1(n377), .B2(n354), .ZN(n221) );
  OAI21_X1 U476 ( .B1(n251), .B2(n386), .A(n326), .ZN(n214) );
  LOGIC0_X1 U478 ( .Z(n18) );
  NAND2_X2 U479 ( .A1(n184), .A2(n171), .ZN(n290) );
  NOR2_X2 U480 ( .A1(d_internal__acc[35]), .A2(n414), .ZN(n289) );
  NAND2_X2 U481 ( .A1(n182), .A2(n407), .ZN(n297) );
  INV_X2 U482 ( .A(n301), .ZN(n302) );
  //INV_X1 U483 ( .A(n456), .ZN(A_out_proc[18]) );
  NOR2_X2 U484 ( .A1(d_internal__acc[21]), .A2(n409), .ZN(n306) );
  NOR2_X2 U485 ( .A1(n306), .A2(n305), .ZN(n308) );
  NAND2_X2 U486 ( .A1(n308), .A2(n307), .ZN(n145) );
  //INV_X1 U487 ( .A(n419), .ZN(A_out_proc[24]) );
  //INV_X1 U488 ( .A(n480), .ZN(A_out_proc[12]) );
  //INV_X1 U489 ( .A(n479), .ZN(A_out_proc[19]) );
  //INV_X1 U490 ( .A(n424), .ZN(A_out_proc[1]) );
  NOR4_X1 U491 ( .A1(state_out_of_wrapper[1]), .A2(n397), .A3(
        state_out_of_wrapper[2]), .A4(count0[6]), .ZN(n317) );
  NAND4_X1 U492 ( .A1(count0[0]), .A2(count0[4]), .A3(count0[1]), .A4(
        count0[5]), .ZN(n313) );
  NOR4_X1 U493 ( .A1(count0[8]), .A2(count0[7]), .A3(n314), .A4(n313), .ZN(
        n316) );
  AOI22_X1 U494 ( .A1(n351), .A2(B_in_to_wrapper[11]), .B1(B_in_to_wrapper[12]), .B2(n350), .ZN(n324) );
  OAI21_X1 U495 ( .B1(n247), .B2(n386), .A(n324), .ZN(n216) );
  //INV_X1 U496 ( .A(n488), .ZN(A_out_proc[3]) );
  INV_X1 U497 ( .A(B_in_to_wrapper[3]), .ZN(n371) );
  INV_X1 U498 ( .A(B_in_to_wrapper[0]), .ZN(n368) );
  INV_X1 U499 ( .A(A_in_to_wrapper[5]), .ZN(n353) );
  INV_X1 U500 ( .A(A_in_to_wrapper[3]), .ZN(n380) );
  INV_X1 U501 ( .A(A_in_to_wrapper[2]), .ZN(n354) );
  INV_X1 U502 ( .A(A_in_to_wrapper[1]), .ZN(n355) );
  INV_X1 U503 ( .A(A_in_to_wrapper[4]), .ZN(n382) );
  INV_X1 U504 ( .A(A_in_to_wrapper[0]), .ZN(n356) );
  INV_X1 U505 ( .A(A_in_to_wrapper[7]), .ZN(n389) );
  //INV_X1 U506 ( .A(n487), .ZN(A_out_proc[4]) );
  //INV_X1 U507 ( .A(n486), .ZN(A_out_proc[5]) );
  //INV_X1 U508 ( .A(n484), .ZN(A_out_proc[6]) );
  //INV_X1 U509 ( .A(n483), .ZN(A_out_proc[7]) );
  //INV_X1 U510 ( .A(n474), .ZN(A_out_proc[8]) );
  //INV_X1 U511 ( .A(n471), .ZN(A_out_proc[9]) );
  //INV_X1 U512 ( .A(n448), .ZN(A_out_proc[14]) );
  //INV_X1 U513 ( .A(n421), .ZN(A_out_proc[17]) );
  //INV_X1 U514 ( .A(n489), .ZN(A_out_proc[13]) );
  //INV_X1 U515 ( .A(n473), .ZN(A_out_proc[15]) );
  NAND2_X2 U516 ( .A1(n361), .A2(n360), .ZN(n442) );
  INV_X4 U517 ( .A(n449), .ZN(A_out[25]) );
  INV_X4 U518 ( .A(n430), .ZN(n138) );
  INV_X4 U519 ( .A(n466), .ZN(n151) );
  INV_X4 U520 ( .A(n426), .ZN(n141) );
  INV_X4 U521 ( .A(n429), .ZN(n133) );
  INV_X4 U522 ( .A(n428), .ZN(n144) );
  INV_X4 U523 ( .A(n427), .ZN(n128) );
  INV_X4 U524 ( .A(n403), .ZN(n139) );
  INV_X4 U525 ( .A(n425), .ZN(n129) );
  INV_X4 U526 ( .A(n388), .ZN(B_out[14]) );
  INV_X4 U527 ( .A(n406), .ZN(n124) );
  INV_X4 U528 ( .A(n453), .ZN(A_out[10]) );
  INV_X4 U529 ( .A(n460), .ZN(A_out[8]) );
  INV_X4 U530 ( .A(n434), .ZN(n136) );
  INV_X4 U531 ( .A(n499), .ZN(A_out[1]) );
  INV_X4 U532 ( .A(n423), .ZN(n142) );
  OAI222_X1 U533 ( .A1(n377), .A2(n369), .B1(n386), .B2(n437), .C1(n376), .C2(
        n368), .ZN(n205) );
  INV_X1 U534 ( .A(B_in_to_wrapper[2]), .ZN(n370) );
  OAI222_X1 U535 ( .A1(n370), .A2(n377), .B1(n386), .B2(n196), .C1(n376), .C2(
        n369), .ZN(n206) );
  OAI222_X1 U536 ( .A1(n371), .A2(n377), .B1(n386), .B2(n248), .C1(n376), .C2(
        n370), .ZN(n207) );
  INV_X1 U537 ( .A(B_in_to_wrapper[5]), .ZN(n374) );
  INV_X1 U538 ( .A(B_out[5]), .ZN(n373) );
  INV_X1 U539 ( .A(B_in_to_wrapper[4]), .ZN(n372) );
  OAI222_X1 U540 ( .A1(n374), .A2(n377), .B1(n386), .B2(n373), .C1(n376), .C2(
        n372), .ZN(n209) );
  INV_X1 U541 ( .A(B_in_to_wrapper[6]), .ZN(n375) );
  OAI222_X1 U542 ( .A1(n375), .A2(n377), .B1(n386), .B2(n438), .C1(n376), .C2(
        n374), .ZN(n210) );
  INV_X1 U543 ( .A(B_in_to_wrapper[7]), .ZN(n378) );
  OAI222_X1 U544 ( .A1(n378), .A2(n377), .B1(n386), .B2(n250), .C1(n376), .C2(
        n375), .ZN(n211) );
  INV_X1 U545 ( .A(A_in_to_wrapper[11]), .ZN(n381) );
  OAI222_X1 U546 ( .A1(n381), .A2(n390), .B1(n380), .B2(n387), .C1(n386), .C2(
        n435), .ZN(n230) );
  INV_X1 U547 ( .A(A_in_to_wrapper[12]), .ZN(n383) );
  OAI222_X1 U548 ( .A1(n383), .A2(n390), .B1(n382), .B2(n387), .C1(n386), .C2(
        n425), .ZN(n231) );
  INV_X1 U549 ( .A(A_in_to_wrapper[14]), .ZN(n385) );
  OAI222_X1 U550 ( .A1(n385), .A2(n390), .B1(n384), .B2(n387), .C1(n386), .C2(
        n478), .ZN(n233) );
  INV_X1 U551 ( .A(A_in_to_wrapper[15]), .ZN(n393) );
  OAI222_X1 U552 ( .A1(n393), .A2(n390), .B1(n389), .B2(n387), .C1(n386), .C2(
        n464), .ZN(n234) );
  INV_X2 U241 ( .A(n404), .ZN(n273) );
  DFFR_X1 \c_reg_reg[0]  ( .D(n255), .CK(clk), .RN(net23470), .QN(P[0]), .Q()
         );
  DFFR_X1 \c_reg_reg[1]  ( .D(n256), .CK(clk), .RN(net23470), .QN(P[1]), .Q()
         );
  INV_X2 U268 ( .A(n287), .ZN(n288) );
  INV_X1 U240 ( .A(d_internal__acc_13), .ZN(n359) );
  INV_X1 U251 ( .A(n387), .ZN(n351) );
  BUF_X1 U264 ( .A(n392), .Z(n175) );
  NAND2_X1 U265 ( .A1(d_internal__acc[23]), .A2(n407), .ZN(n269) );
  AOI21_X1 U267 ( .B1(n317), .B2(n316), .A(n315), .ZN(n387) );
  OR2_X1 U278 ( .A1(d_internal__acc_8), .A2(n414), .ZN(n255) );
  OR2_X1 U294 ( .A1(d_internal__acc_10), .A2(n414), .ZN(n270) );
  LOGIC1_X1 U309 ( .Z(net23470) );
  INV_X4 U367 ( .A(d_internal__acc[30]), .ZN(n184) );
  /* 
  dummy_load my_dummy ( .A_out({n501, A_out[24:19], n505, A_out[17:14], n508, 
        A_out[12:11], n509, n510, n511, n18, n18, n18, n18, n18, n18, n18, n18}), .B_out({n412, n477, B_out[12:8], n18, n18, n18, n18, n18, n18, n18, n18}), 
        .\A_out_proc[23]_BAR (n401), .\A_out_proc[0] (A_out_proc[0]), 
        .\A_out_proc[20] (A_out_proc[20]), .\A_out_proc[10] (A_out_proc[10]), 
        .\A_out_proc[11] (A_out_proc[11]), .\A_out_proc[24]_BAR (n419), 
        .\A_out_proc[17]_BAR (n421), .\A_out_proc[1]_BAR (n424), 
        .\A_out_proc[14]_BAR (n448), .\A_out_proc[18]_BAR (n456), 
        .\A_out_proc[16] (A_out_proc[16]), .\A_out_proc[19]_BAR (n479), 
        .\A_out_proc[12]_BAR (n480), .\A_out_proc[7]_BAR (n483), 
        .\A_out_proc[6]_BAR (n484), .\A_out_proc[5]_BAR (n486), 
        .\A_out_proc[4]_BAR (n487), .\A_out_proc[3]_BAR (n488), 
        .\A_out_proc[15]_BAR (n473), .\A_out_proc[9]_BAR (n471), 
        .\A_out_proc[8]_BAR (n474), .\A_out_proc[21] (A_out_proc[21]), 
        .\A_out_proc[2] (A_out_proc[2]), .\A_out_proc[13]_BAR (n489), 
        .\A_out_proc[22] (n445) );
   */
   conf_int_mul__noFF__arch_agnos_OP_BITWIDTH18_DATA_PATH_BITWIDTH26__acc mul__inst ( 
        .clk(clk), .racc(n18), .rapx(n18), .a({A_out[25], n138, n151, n141, 
        n133, n144, n128, A_out[18], n134, n121, n120, n122, A_out[13], n129, 
        n131, A_out[10:0]}), .b({B_out[14:13], n139, n148, n124, n149, n482, 
        n150, B_out[6], n142, n485, n136, B_out[2:0]}), .\d[40] (), .\d[39] (
        d_internal__acc[39]), .\d[36] (d_internal__acc[36]), .\d[34] (
        d_internal__acc[34]), .\d[32] (d_internal__acc[32]), .\d[29] (
        d_internal__acc[29]), .\d[25] (d_internal__acc[25]), .\d[23] (
        d_internal__acc[23]), .\d[11] (d_internal__acc_11), .\d[7] (), 
        .\d[6] (), .\d[5] (), .\d[4] (), .\d[3] (), .\d[2] (), .\d[1] (), 
        .\d[0] (), .\d[37]_BAR (d_internal__acc[37]), .\d[30]_BAR (
        d_internal__acc[30]), .\d[24]_BAR (d_internal__acc[24]), .\d[21]_BAR (
        d_internal__acc[21]), .\d[20]_BAR (d_internal__acc[20]), .\d[14]_BAR (
        d_internal__acc_14), .\d[9]_BAR (d_internal__acc_9), .\d[8]_BAR (
        d_internal__acc_8), .\d[28] (d_internal__acc[28]), .\d[27]_BAR (
        d_internal__acc[27]), .\d[31]_BAR (d_internal__acc[31]), .\d[17] (
        d_internal__acc_17), .\d[13]_BAR (d_internal__acc_13), .\d[35]_BAR (
        d_internal__acc[35]), .\d[19] (n164), .\d[22]_BAR (d_internal__acc[22]), .\d[15]_BAR (n417), .\d[18] (d_internal__acc_18), .\d[10]_BAR (
        d_internal__acc_10), .\d[16]_BAR (d_internal__acc_16), .\d[33] (
        d_internal__acc[33]), .\d[38]_BAR (d_internal__acc[38]), .\d[12]_BAR (
        d_internal__acc_12), .\d[26] (d_internal__acc[26]) );
  DFFR_X1 \a_reg_reg[2]  ( .D(n221), .CK(clk), .RN(n444), .QN(n431), .Q(
        A_out[2]) );
  NAND2_X1 U274 ( .A1(n463), .A2(rapx), .ZN(n327) );
  NAND2_X1 U280 ( .A1(d_internal__acc_11), .A2(n171), .ZN(n198) );
  NAND2_X1 U289 ( .A1(n322), .A2(n321), .ZN(n390) );
  INV_X1 U356 ( .A(n443), .ZN(B_out[0]) );
  INV_X1 U242 ( .A(n357), .ZN(n330) );
  NAND2_X1 U244 ( .A1(n390), .A2(n387), .ZN(n357) );
  INV_X1 U249 ( .A(rstP), .ZN(n284) );
  OR2_X1 U254 ( .A1(acc__sel), .A2(rstP), .ZN(n286) );
  INV_X1 U255 ( .A(n490), .ZN(n322) );
  OAI21_X1 U270 ( .B1(state_out_of_wrapper[2]), .B2(state_out_of_wrapper[1]), 
        .A(n318), .ZN(n490) );
endmodule


module conf_int_mul__noFF__arch_agnos ( clk, racc, rapx, a, b, d);
   parameter OP_BITWIDTH = 16; 
   parameter DATA_PATH_BITWIDTH = 24;
   
   input clk;
   input racc;
   input rapx;
   input [DATA_PATH_BITWIDTH -1: 0] a;
   input [DATA_PATH_BITWIDTH -1 - 11: 0] b;
   //output [(DATA_PATH_BITWIDTH + DATA_PATH_BITWIDTH ) - 1 - 11 : 0] d;
   output [(DATA_PATH_BITWIDTH - 8+ DATA_PATH_BITWIDTH - 8) - 1 - 11 : 0] d;
   assign d = $signed(a[25:8]) * $signed(b[14:8]);
endmodule


module conf_int_mul__noFF__arch_agnos__w_wrapper(A_in_to_wrapper, B_in_to_wrapper, state_in_to_wrapper, rstP, clk, racc,rapx, P, count0, state_out_of_wrapper, acc__sel);
   parameter OP_BITWIDTH = 16; //operator bit width
   parameter DATA_PATH_BITWIDTH = 24; //flip flop Bit width
   
   input [DATA_PATH_BITWIDTH -1: 0] A_in_to_wrapper;
   input [DATA_PATH_BITWIDTH -1 - 11: 0] B_in_to_wrapper;
   input [8:0] count0;
   input [2:0] state_in_to_wrapper;      
   output [2:0] state_out_of_wrapper;      
   input acc__sel;
   wire [(DATA_PATH_BITWIDTH - 8 + DATA_PATH_BITWIDTH - 8) - 1 -11:0] d_internal__apx;
   input rstP; 
   input clk;
   input racc; //accurate bits reset  
   input rapx; //apx bits reset
   output [31:0] P; 
   wire [DATA_PATH_BITWIDTH -1: 0] A_out;
   wire [DATA_PATH_BITWIDTH -1 - 11: 0] B_out;

//wire [DATA_PATH_BITWIDTH:0] d__acc;
// synopsys dc_script_begin
 //set_dont_touch mul__inst__acc
 // synopsys dc_script_end
conf_int_mul__noFF__arch_agnos #(OP_BITWIDTH, DATA_PATH_BITWIDTH) mul__inst__apx(.clk(clk), .racc(racc), .rapx(rapx),.a(A_out), .b(B_out), .d(d_internal__apx));



//conf_int_mul__noFF__arch_agnos__w_wrapper #(OP_BITWIDTH, DATA_PATH_BITWIDTH) mul__inst__acc(A_in_to_wrapper, B_in_to_wrapper, state_in_to_wrapper, rstP, clk, racc,rapx, P, count0, state_out_of_wrapper, d_internal__apx, acc__sel, A_out, B_out);
conf_int_mul__noFF__arch_agnos__w_wrapper_OP_BITWIDTH18_DATA_PATH_BITWIDTH26__acc mul__inst__acc( 
        A_in_to_wrapper, B_in_to_wrapper, state_in_to_wrapper, rstP, clk, racc, 
        rapx, P, count0, state_out_of_wrapper, d_internal__apx, acc__sel, 
        A_out, B_out);



//--- for testing purposes
//--- duplicate
//assign d = d__ignore;
/*
// ---- non duplicates
//--- F:DN acc
//assign d = a*b; 

//-- F:DN apx
assign d[63:16] = a[23:8]*b[23:8]; //apx
assign d[15:0] = 16'b0;
*/

endmodule 
