library verilog;
use verilog.vl_types.all;
entity LOGIC1_X1_func is
    port(
        Z               : out    vl_logic
    );
end LOGIC1_X1_func;
