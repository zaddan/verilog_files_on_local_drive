library verilog;
use verilog.vl_types.all;
entity LOGIC0_X1 is
    port(
        Z               : out    vl_logic
    );
end LOGIC0_X1;
