library verilog;
use verilog.vl_types.all;
entity CLKGATETST_X1_func is
    port(
        CK              : in     vl_logic;
        E               : in     vl_logic;
        SE              : in     vl_logic;
        GCK             : out    vl_logic
    );
end CLKGATETST_X1_func;
