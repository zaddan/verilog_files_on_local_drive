library verilog;
use verilog.vl_types.all;
entity \conf_int_mul__noFF__arch_agnos_OP_BITWIDTH18_DATA_PATH_BITWIDTH26\ is
    port(
        clk             : in     vl_logic;
        racc            : in     vl_logic;
        rapx            : in     vl_logic;
        a               : in     vl_logic_vector(25 downto 0);
        b               : in     vl_logic_vector(14 downto 0);
        \d_40_\         : out    vl_logic;
        \d_39_\         : out    vl_logic;
        \d_38_\         : out    vl_logic;
        \d_37_\         : out    vl_logic;
        \d_35__BAR\     : out    vl_logic;
        \d_34_\         : out    vl_logic;
        \d_32_\         : out    vl_logic;
        \d_27_\         : out    vl_logic;
        \d_20_\         : out    vl_logic;
        \d_15_\         : out    vl_logic;
        \d_7_\          : out    vl_logic;
        \d_6_\          : out    vl_logic;
        \d_5_\          : out    vl_logic;
        \d_4_\          : out    vl_logic;
        \d_3_\          : out    vl_logic;
        \d_2_\          : out    vl_logic;
        \d_1_\          : out    vl_logic;
        \d_0_\          : out    vl_logic;
        \d_33__BAR\     : out    vl_logic;
        \d_30__BAR\     : out    vl_logic;
        \d_9_\          : out    vl_logic;
        \d_31__BAR\     : out    vl_logic;
        \d_28__BAR\     : out    vl_logic;
        \d_25__BAR\     : out    vl_logic;
        \d_11__BAR\     : out    vl_logic;
        \d_36_\         : out    vl_logic;
        \d_26__BAR\     : out    vl_logic;
        \d_19_\         : out    vl_logic;
        \d_29__BAR\     : out    vl_logic;
        \d_18__BAR\     : out    vl_logic;
        \d_10__BAR\     : out    vl_logic;
        \d_24_\         : out    vl_logic;
        \d_8_\          : out    vl_logic;
        \d_13__BAR\     : out    vl_logic;
        \d_17_\         : out    vl_logic;
        \d_16_\         : out    vl_logic;
        \d_22_\         : out    vl_logic;
        \d_14__BAR\     : out    vl_logic;
        \d_23_\         : out    vl_logic;
        \d_21__BAR\     : out    vl_logic;
        \d_12__BAR\     : out    vl_logic
    );
end \conf_int_mul__noFF__arch_agnos_OP_BITWIDTH18_DATA_PATH_BITWIDTH26\;
